@comment $OpenBSD: PLIST.sv,v 1.2 2002/04/15 06:53:53 espie Exp $
share/apps/ktuberling/sounds/sv/brosch.wav
share/apps/ktuberling/sounds/sv/cigarr.wav
share/apps/ktuberling/sounds/sv/fluga.wav
share/apps/ktuberling/sounds/sv/glasogon.wav
share/apps/ktuberling/sounds/sv/halsband.wav
share/apps/ktuberling/sounds/sv/halsduk.wav
share/apps/ktuberling/sounds/sv/har.wav
share/apps/ktuberling/sounds/sv/hatt.wav
share/apps/ktuberling/sounds/sv/horn.wav
share/apps/ktuberling/sounds/sv/klocka.wav
share/apps/ktuberling/sounds/sv/mun.wav
share/apps/ktuberling/sounds/sv/mustasch.wav
share/apps/ktuberling/sounds/sv/nasa.wav
share/apps/ktuberling/sounds/sv/oga.wav
share/apps/ktuberling/sounds/sv/ogonbryn.wav
share/apps/ktuberling/sounds/sv/ora.wav
share/apps/ktuberling/sounds/sv/orhange.wav
share/apps/ktuberling/sounds/sv/pingvin.wav
share/apps/ktuberling/sounds/sv/potatismannen.wav
share/apps/ktuberling/sounds/sv/rosett.wav
share/apps/ktuberling/sounds/sv/slips.wav
share/apps/ktuberling/sounds/sv/solglasogon.wav
${DOC}KRegExpEditor/altntool.png
${DOC}KRegExpEditor/anychartool.png
${DOC}KRegExpEditor/boundarytools.png
${DOC}KRegExpEditor/charactertool.png
${DOC}KRegExpEditor/common
${DOC}KRegExpEditor/compoundtool.png
${DOC}KRegExpEditor/${C}
${DOC}KRegExpEditor/${I}
${DOC}KRegExpEditor/linestartendtool.png
${DOC}KRegExpEditor/lookaheadtools.png
${DOC}KRegExpEditor/repeattool.png
${DOC}KRegExpEditor/theEditor.png
${DOC}aktion/common
${DOC}aktion/${C}
${DOC}aktion/${I}
${DOC}amor/common
${DOC}amor/${C}
${DOC}amor/${I}
${DOC}ark/common
${DOC}ark/${C}
${DOC}ark/${I}
${DOC}artsbuilder/apis.docbook
${DOC}artsbuilder/arts-structure.png
${DOC}artsbuilder/artsbuilder.docbook
${DOC}artsbuilder/common
${DOC}artsbuilder/detail.docbook
${DOC}artsbuilder/digitalaudio.docbook
${DOC}artsbuilder/faq.docbook
${DOC}artsbuilder/future.docbook
${DOC}artsbuilder/glossary.docbook
${DOC}artsbuilder/gui.docbook
${DOC}artsbuilder/helping.docbook
${DOC}artsbuilder/images/Synth_AMAN_PLAY.png
${DOC}artsbuilder/images/Synth_AMAN_RECORD.png
${DOC}artsbuilder/images/Synth_BRICKWALL_LIMITER.png
${DOC}artsbuilder/images/Synth_CAPTURE.png
${DOC}artsbuilder/images/Synth_DATA.png
${DOC}artsbuilder/images/Synth_FREEVERB.png
${DOC}artsbuilder/images/Synth_FX_CFLANGER.png
${DOC}artsbuilder/images/Synth_MIDI_TEST.png
${DOC}artsbuilder/images/Synth_MOOG_VCF.png
${DOC}artsbuilder/images/Synth_MULTI_ADD.png
${DOC}artsbuilder/images/Synth_NOISE.png
${DOC}artsbuilder/images/Synth_PITCH_SHIFT.png
${DOC}artsbuilder/images/Synth_RECORD.png
${DOC}artsbuilder/images/Synth_TREMOLO.png
${DOC}artsbuilder/images/Synth_WAVE_PULSE.png
${DOC}artsbuilder/images/Synth_WAVE_SOFTSAW.png
${DOC}artsbuilder/${C}
${DOC}artsbuilder/${I}
${DOC}artsbuilder/mcop.docbook
${DOC}artsbuilder/midi.docbook
${DOC}artsbuilder/midiintro.docbook
${DOC}artsbuilder/modules.docbook
${DOC}artsbuilder/porting.docbook
${DOC}artsbuilder/references.docbook
${DOC}artsbuilder/tools.docbook
${DOC}cervisia/checkout.png
${DOC}cervisia/commit.png
${DOC}cervisia/common
${DOC}cervisia/diff.png
${DOC}cervisia/history.png
${DOC}cervisia/import.png
${DOC}cervisia/${C}
${DOC}cervisia/${I}
${DOC}cervisia/logtree.png
${DOC}cervisia/mainview.png
${DOC}cervisia/resolve.png
${DOC}cervisia/updatetag.png
${DOC}common/1.png
${DOC}common/10.png
${DOC}common/2.png
${DOC}common/3.png
${DOC}common/4.png
${DOC}common/5.png
${DOC}common/6.png
${DOC}common/7.png
${DOC}common/8.png
${DOC}common/9.png
${DOC}common/artistic-license.html
${DOC}common/bottom1.png
${DOC}common/bottom2.png
${DOC}common/bsd-license.html
${DOC}common/doctop1.png
${DOC}common/doctop1a.png
${DOC}common/doctop1b.png
${DOC}common/doctop2.png
${DOC}common/fdl-license
${DOC}common/fdl-license.html
${DOC}common/fdl-translated.html
${DOC}common/gpl-license
${DOC}common/gpl-license.html
${DOC}common/gpl-translated.html
${DOC}common/kde-common.css
${DOC}common/kde-default.css
${DOC}common/kde-localised.css
${DOC}common/kde-localised.css.template
${DOC}common/kde-web.css
${DOC}common/lgpl-license
${DOC}common/lgpl-license.html
${DOC}common/lgpl-translated.html
${DOC}common/logotp3.png
${DOC}common/qpl-license.html
${DOC}common/shadow.png
${DOC}common/web-docbottom.png
${DOC}common/web-doctop.png
${DOC}common/x11-license.html
${DOC}common/xml.dcl
${DOC}kab/common
${DOC}kab/${C}
${DOC}kab/${I}
${DOC}kab/kab-edit.png
${DOC}kab/kab-using.png
${DOC}kaddressbook/common
${DOC}kaddressbook/${C}
${DOC}kaddressbook/${I}
${DOC}kalarm/alarmmessage.png
${DOC}kalarm/common
${DOC}kalarm/editwindow.png
${DOC}kalarm/${C}
${DOC}kalarm/${I}
${DOC}kalarm/mainwindow.png
${DOC}kandy/common
${DOC}kandy/${C}
${DOC}kandy/${I}
${DOC}karm/common
${DOC}karm/${C}
${DOC}karm/${I}
${DOC}kasteroids/common
${DOC}kasteroids/${C}
${DOC}kasteroids/${I}
${DOC}kate-plugins/common
${DOC}kate-plugins/helloworld.docbook
${DOC}kate-plugins/htmltools.docbook
${DOC}kate-plugins/${C}
${DOC}kate-plugins/${I}
${DOC}kate-plugins/insertcommand.docbook
${DOC}kate-plugins/openheader.docbook
${DOC}kate-plugins/projectmanager.docbook
${DOC}kate-plugins/textfilter.docbook
${DOC}kate-plugins/xmltools.docbook
${DOC}kate/advanced.docbook
${DOC}kate/common
${DOC}kate/configdialog01.png
${DOC}kate/configdialog02.png
${DOC}kate/configuring.docbook
${DOC}kate/fundamentals.docbook
${DOC}kate/highlighting.docbook
${DOC}kate/${C}
${DOC}kate/${I}
${DOC}kate/kate.png
${DOC}kate/mdi.docbook
${DOC}kate/menus.docbook
${DOC}kate/mimetypechooser.png
${DOC}kate/part.docbook
${DOC}kate/plugins.docbook
${DOC}kate/regular-expressions.docbook
${DOC}katomic/common
${DOC}katomic/${C}
${DOC}katomic/${I}
${DOC}kbabel/common
${DOC}kbabel/${C}
${DOC}kbabel/${I}
${DOC}kbabel/snap1.png
${DOC}kbabel/snap_catalogmanager.png
${DOC}kbackgammon/common
${DOC}kbackgammon/${C}
${DOC}kbackgammon/${I}
${DOC}kbattleship/common
${DOC}kbattleship/${C}
${DOC}kbattleship/${I}
${DOC}kblackbox/common
${DOC}kblackbox/${C}
${DOC}kblackbox/${I}
${DOC}kbounce/common
${DOC}kbounce/${C}
${DOC}kbounce/${I}
${DOC}kcalc/common
${DOC}kcalc/${C}
${DOC}kcalc/${I}
${DOC}kcoloredit/common
${DOC}kcoloredit/${C}
${DOC}kcoloredit/${I}
${DOC}kcontrol/common
${DOC}kcontrol/${C}
${DOC}kcontrol/${I}
${DOC}kcontrol/kalarmd.docbook
${DOC}kcontrol/kcmaccess.docbook
${DOC}kcontrol/kcmaction.docbook
${DOC}kcontrol/kcmbackgnd.docbook
${DOC}kcontrol/kcmbatmon.docbook
${DOC}kcontrol/kcmbell.docbook
${DOC}kcontrol/kcmblockdev.docbook
${DOC}kcontrol/kcmcache.docbook
${DOC}kcontrol/kcmcolor.docbook
${DOC}kcontrol/kcmcookie.docbook
${DOC}kcontrol/kcmcrypto.docbook
${DOC}kcontrol/kcmcss.docbook
${DOC}kcontrol/kcmdatetime.docbook
${DOC}kcontrol/kcmdesktop.docbook
${DOC}kcontrol/kcmdeviceinfo.docbook
${DOC}kcontrol/kcmdmainfo.docbook
${DOC}kcontrol/kcmebrowse.docbook
${DOC}kcontrol/kcmemail.docbook
${DOC}kcontrol/kcmenergy.docbook
${DOC}kcontrol/kcmfile.docbook
${DOC}kcontrol/kcmfileman.docbook
${DOC}kcontrol/kcmfontinst.docbook
${DOC}kcontrol/kcmfonts.docbook
${DOC}kcontrol/kcmhelp${I}
${DOC}kcontrol/kcmicon.docbook
${DOC}kcontrol/kcmintinfo.docbook
${DOC}kcontrol/kcmioportinfo.docbook
${DOC}kcontrol/kcmkbd.docbook
${DOC}kcontrol/kcmkbrowse.docbook
${DOC}kcontrol/kcmkeybind.docbook
${DOC}kcontrol/kcmkonsole.docbook
${DOC}kcontrol/kcmkwintheme.docbook
${DOC}kcontrol/kcmlaunch.docbook
${DOC}kcontrol/kcmlisa.docbook
${DOC}kcontrol/kcmlocate.docbook
${DOC}kcontrol/kcmloginmanage.docbook
${DOC}kcontrol/kcmlowbatcrit.docbook
${DOC}kcontrol/kcmlowbatwarn.docbook
${DOC}kcontrol/kcmmemoryinfo.docbook
${DOC}kcontrol/kcmmidi.docbook
${DOC}kcontrol/kcmmixer.docbook
${DOC}kcontrol/kcmmouse.docbook
${DOC}kcontrol/kcmnetscapeplugins.docbook
${DOC}kcontrol/kcmnics.docbook
${DOC}kcontrol/kcmpanel.docbook
${DOC}kcontrol/kcmpartitioninfo.docbook
${DOC}kcontrol/kcmpasswd.docbook
${DOC}kcontrol/kcmpciinfo.docbook
${DOC}kcontrol/kcmpcmcia.docbook
${DOC}kcontrol/kcmpowerctrl.docbook
${DOC}kcontrol/kcmprocinfo.docbook
${DOC}kcontrol/kcmproxie.docbook
${DOC}kcontrol/kcmscnsave.docbook
${DOC}kcontrol/kcmscsiinfo.docbook
${DOC}kcontrol/kcmsessionman.docbook
${DOC}kcontrol/kcmsmbstat.docbook
${DOC}kcontrol/kcmsndinfo.docbook
${DOC}kcontrol/kcmsndsrv.docbook
${DOC}kcontrol/kcmsocks.docbook
${DOC}kcontrol/kcmspellchecking.docbook
${DOC}kcontrol/kcmstyle.docbook
${DOC}kcontrol/kcmsysnotify.docbook
${DOC}kcontrol/kcmtalk.docbook
${DOC}kcontrol/kcmtaskbar.docbook
${DOC}kcontrol/kcmusb.docbook
${DOC}kcontrol/kcmuseragent.docbook
${DOC}kcontrol/kcmwinshare.docbook
${DOC}kcontrol/kcmxmlrpc.docbook
${DOC}kcontrol/kcmxservinfo.docbook
${DOC}kcontrol/nettimeouts.docbook
${DOC}kcontrol/printmanager.docbook
${DOC}kcontrol/printsystem.docbook
${DOC}kcontrol/protocols.docbook
${DOC}kcontrol/screenshot.png
${DOC}kcontrol/systemcontrol.docbook
${DOC}kcontrol/thememgr.docbook
${DOC}kcron/common
${DOC}kcron/${C}
${DOC}kcron/${I}
${DOC}kcron/kcron.png
${DOC}kcron/kcronstart.png
${DOC}kcron/newtask.png
${DOC}kcron/newvariable.png
${DOC}kcron/print.png
${DOC}kdat/common
${DOC}kdat/${C}
${DOC}kdat/${I}
${DOC}kdebugdialog/common
${DOC}kdebugdialog/${C}
${DOC}kdebugdialog/${I}
${DOC}kdeprint/add-printer-wiz.docbook
${DOC}kdeprint/common
${DOC}kdeprint/cups-config.docbook
${DOC}kdeprint/cups-filterarchitecture-kivio-70Percent-scaled.png
${DOC}kdeprint/cupsaddprinterwizard1.png
${DOC}kdeprint/cupsaddprinterwizard2_backendselection.png
${DOC}kdeprint/cupsoptions.docbook
${DOC}kdeprint/extensions.docbook
${DOC}kdeprint/external-command.docbook
${DOC}kdeprint/final-word.docbook
${DOC}kdeprint/getting-started.docbook
${DOC}kdeprint/highlights.docbook
${DOC}kdeprint/${C}
${DOC}kdeprint/${I}
${DOC}kdeprint/kprinter-kivio.png
${DOC}kdeprint/kprinter_called_from_run_command.png
${DOC}kdeprint/lpd.docbook
${DOC}kdeprint/lpr-bsd.docbook
${DOC}kdeprint/lprng.docbook
${DOC}kdeprint/rlpr.docbook
${DOC}kdeprint/tech-overview.docbook
${DOC}kdeprint/theory.docbook
${DOC}kdesu/common
${DOC}kdesu/${C}
${DOC}kdesu/${I}
${DOC}kdevelop/tip.database
${DOC}kdf/common
${DOC}kdf/${C}
${DOC}kdf/${I}
${DOC}kdf/kdf.png
${DOC}kdf/kdf_config.png
${DOC}kdict/applet.png
${DOC}kdict/common
${DOC}kdict/conf.png
${DOC}kdict/${C}
${DOC}kdict/${I}
${DOC}kdict/mainwin.png
${DOC}kdict/seteditor.png
${DOC}kdm/common
${DOC}kdm/${C}
${DOC}kdm/${I}
${DOC}kdvi/common
${DOC}kdvi/${C}
${DOC}kdvi/${I}
${DOC}kdvi/optionrequester1.png
${DOC}kdvi/optionrequester2.png
${DOC}kedit/common
${DOC}kedit/${C}
${DOC}kedit/${I}
${DOC}kenolaba/common
${DOC}kenolaba/${C}
${DOC}kenolaba/${I}
${DOC}kfind/common
${DOC}kfind/${C}
${DOC}kfind/${I}
${DOC}kfloppy/common
${DOC}kfloppy/${C}
${DOC}kfloppy/${I}
${DOC}kformula/common
${DOC}kformula/${C}
${DOC}kformula/${I}
${DOC}kfouleggs/common
${DOC}kfouleggs/${C}
${DOC}kfouleggs/${I}
${DOC}kfract/common
${DOC}kfract/${C}
${DOC}kfract/${I}
${DOC}kgeo/common
${DOC}kgeo/${C}
${DOC}kgeo/${I}
${DOC}kghostview/common
${DOC}kghostview/${C}
${DOC}kghostview/${I}
${DOC}khangman/common
${DOC}khangman/${C}
${DOC}khangman/${I}
${DOC}khelpcenter/common
${DOC}khelpcenter/contact.docbook
${DOC}khelpcenter/faq/about.docbook
${DOC}khelpcenter/faq/common
${DOC}khelpcenter/faq/configkde.docbook
${DOC}khelpcenter/faq/contrib.docbook
${DOC}khelpcenter/faq/desktop.docbook
${DOC}khelpcenter/faq/filemng.docbook
${DOC}khelpcenter/faq/getkde.docbook
${DOC}khelpcenter/faq/${C}
${DOC}khelpcenter/faq/${I}
${DOC}khelpcenter/faq/install.docbook
${DOC}khelpcenter/faq/intro.docbook
${DOC}khelpcenter/faq/kdeapps.docbook
${DOC}khelpcenter/faq/misc.docbook
${DOC}khelpcenter/faq/moreinfo.docbook
${DOC}khelpcenter/faq/nonkdeapps.docbook
${DOC}khelpcenter/faq/notrelated.docbook
${DOC}khelpcenter/faq/panel.docbook
${DOC}khelpcenter/faq/tips.docbook
${DOC}khelpcenter/faq/winmng.docbook
${DOC}khelpcenter/glossary/common
${DOC}khelpcenter/glossary/${C}
${DOC}khelpcenter/glossary/${I}
${DOC}khelpcenter/glossary/kdeprintingglossary.docbook
${DOC}khelpcenter/help.docbook
${DOC}khelpcenter/${C}
${DOC}khelpcenter/${I}
${DOC}khelpcenter/links.docbook
${DOC}khelpcenter/quickstart/common
${DOC}khelpcenter/quickstart/${C}
${DOC}khelpcenter/quickstart/${I}
${DOC}khelpcenter/support.docbook
${DOC}khelpcenter/userguide/about-desktop.docbook
${DOC}khelpcenter/userguide/common
${DOC}khelpcenter/userguide/first-impressions.docbook
${DOC}khelpcenter/userguide/getting-started.docbook
${DOC}khelpcenter/userguide/history.docbook
${DOC}khelpcenter/userguide/${C}
${DOC}khelpcenter/userguide/${I}
${DOC}khelpcenter/userguide/installation.docbook
${DOC}khelpcenter/userguide/intro.docbook
${DOC}khelpcenter/userguide/kdeadmin-apps.docbook
${DOC}khelpcenter/userguide/kdebase-apps.docbook
${DOC}khelpcenter/userguide/kdeedu-apps.docbook
${DOC}khelpcenter/userguide/kdegames-apps.docbook
${DOC}khelpcenter/userguide/kdegraphics-apps.docbook
${DOC}khelpcenter/userguide/kdemultimedia-apps.docbook
${DOC}khelpcenter/userguide/kdenetwork-apps.docbook
${DOC}khelpcenter/userguide/kdepim-apps.docbook
${DOC}khelpcenter/userguide/kdetoys-apps.docbook
${DOC}khelpcenter/userguide/kdeutils-apps.docbook
${DOC}khelpcenter/userguide/koffice-apps.docbook
${DOC}khelpcenter/userguide/more-help.docbook
${DOC}khelpcenter/userguide/shortcuts.docbook
${DOC}khelpcenter/userguide/staff.docbook
${DOC}khelpcenter/userguide/ug-faq.docbook
${DOC}khelpcenter/visualdict/common
${DOC}khelpcenter/visualdict/${C}
${DOC}khelpcenter/visualdict/${I}
${DOC}khelpcenter/welcome.docbook
${DOC}khelpcenter/whatiskde.docbook
${DOC}khexedit/common
${DOC}khexedit/${C}
${DOC}khexedit/${I}
${DOC}khexedit/khexedit1.png
${DOC}kicker-applets/common
${DOC}kicker-applets/${C}
${DOC}kicker-applets/${I}
${DOC}kicker-applets/kolourpicker.docbook
${DOC}kicker-applets/ktimemon.docbook
${DOC}kicker/common
${DOC}kicker/${C}
${DOC}kicker/${I}
${DOC}kiconedit/common
${DOC}kiconedit/${C}
${DOC}kiconedit/${I}
${DOC}kioslave/audiocd.docbook
${DOC}kioslave/bzip.docbook
${DOC}kioslave/bzip2.docbook
${DOC}kioslave/common
${DOC}kioslave/file.docbook
${DOC}kioslave/finger.docbook
${DOC}kioslave/floppy.docbook
${DOC}kioslave/ftp.docbook
${DOC}kioslave/gopher.docbook
${DOC}kioslave/gzip.docbook
${DOC}kioslave/help.docbook
${DOC}kioslave/http.docbook
${DOC}kioslave/https.docbook
${DOC}kioslave/imap.docbook
${DOC}kioslave/imaps.docbook
${DOC}kioslave/${C}
${DOC}kioslave/${I}
${DOC}kioslave/info.docbook
${DOC}kioslave/lan.docbook
${DOC}kioslave/ldap.docbook
${DOC}kioslave/mailto.docbook
${DOC}kioslave/man.docbook
${DOC}kioslave/news.docbook
${DOC}kioslave/nfs.docbook
${DOC}kioslave/nntp.docbook
${DOC}kioslave/pop3.docbook
${DOC}kioslave/pop3s.docbook
${DOC}kioslave/print.docbook
${DOC}kioslave/rdate.docbook
${DOC}kioslave/rlan.docbook
${DOC}kioslave/rlogin.docbook
${DOC}kioslave/sftp.docbook
${DOC}kioslave/smb.docbook
${DOC}kioslave/smtp.docbook
${DOC}kioslave/tar.docbook
${DOC}kioslave/telnet.docbook
${DOC}kioslave/thumbnail.docbook
${DOC}kioslave/webdav.docbook
${DOC}kioslave/webdavs.docbook
${DOC}kit/common
${DOC}kit/${C}
${DOC}kit/${I}
${DOC}kjots/common
${DOC}kjots/${C}
${DOC}kjots/${I}
${DOC}kjumpingcube/common
${DOC}kjumpingcube/${C}
${DOC}kjumpingcube/${I}
${DOC}klettres/common
${DOC}klettres/${C}
${DOC}klettres/${I}
${DOC}klettres/klettres1.png
${DOC}klettres/klettres3.png
${DOC}klines/common
${DOC}klines/${C}
${DOC}klines/${I}
${DOC}klipper/common
${DOC}klipper/${C}
${DOC}klipper/${I}
${DOC}kljettool/common
${DOC}kljettool/${C}
${DOC}kljettool/${I}
${DOC}kljettool/screenshot.png
${DOC}klpq/common
${DOC}klpq/${C}
${DOC}klpq/${I}
${DOC}klprfax/common
${DOC}klprfax/${C}
${DOC}klprfax/${I}
${DOC}kmail/common
${DOC}kmail/${C}
${DOC}kmail/${I}
${DOC}kmenuedit/common
${DOC}kmenuedit/${C}
${DOC}kmenuedit/${I}
${DOC}kmessedwords/common
${DOC}kmessedwords/${C}
${DOC}kmessedwords/${I}
${DOC}kmessedwords/kmw1.png
${DOC}kmessedwords/kmw2.png
${DOC}kmessedwords/kmw3.png
${DOC}kmessedwords/kmw4.png
${DOC}kmid/common
${DOC}kmid/${C}
${DOC}kmid/${I}
${DOC}kmidi/common
${DOC}kmidi/${C}
${DOC}kmidi/${I}
${DOC}kmines/common
${DOC}kmines/${C}
${DOC}kmines/${I}
${DOC}kmines/kmines1.png
${DOC}kmines/kmines2.png
${DOC}kmix/common
${DOC}kmix/${C}
${DOC}kmix/${I}
${DOC}kmoon/common
${DOC}kmoon/${C}
${DOC}kmoon/${I}
${DOC}knewsticker/common
${DOC}knewsticker/contextmenu.png
${DOC}knewsticker/${C}
${DOC}knewsticker/${I}
${DOC}knewsticker/kcmnewsticker-general.png
${DOC}knewsticker/kcmnewsticker-newssources.png
${DOC}knode/common
${DOC}knode/${C}
${DOC}knode/${I}
${DOC}knode/knode-cleanup.png
${DOC}knode/knode-colors-fonts.png
${DOC}knode/knode-composer-attachments.png
${DOC}knode/knode-composer-settings.png
${DOC}knode/knode-edit-filter.png
${DOC}knode/knode-edit-header1.png
${DOC}knode/knode-edit-header2.png
${DOC}knode/knode-filters.png
${DOC}knode/knode-followup.png
${DOC}knode/knode-header-settings.png
${DOC}knode/knode-identity.png
${DOC}knode/knode-mail-account.png
${DOC}knode/knode-new-article.png
${DOC}knode/knode-news-account.png
${DOC}knode/knode-post-settings.png
${DOC}knode/knode-read-news-settings.png
${DOC}knode/knode-reply.png
${DOC}knode/knode-search.png
${DOC}knode/knode-start.png
${DOC}knode/knode-subscribe.png
${DOC}knode/knode-views.png
${DOC}knotes/common
${DOC}knotes/${C}
${DOC}knotes/${I}
${DOC}kodo/common
${DOC}kodo/${C}
${DOC}kodo/${I}
${DOC}koffice/common
${DOC}koffice/${C}
${DOC}koffice/${I}
${DOC}koncd/audiocd.jpg
${DOC}koncd/common
${DOC}koncd/copycd.jpg
${DOC}koncd/imagetype.jpg
${DOC}koncd/${C}
${DOC}koncd/${I}
${DOC}koncd/koncd_logo.jpg
${DOC}koncd/mastercd.jpg
${DOC}koncd/ripcd.jpg
${DOC}koncd/setup.jpg
${DOC}koncd/tools.jpg
${DOC}konq-plugins/archiver.docbook
${DOC}konq-plugins/babel.docbook
${DOC}konq-plugins/common
${DOC}konq-plugins/dirfilter.docbook
${DOC}konq-plugins/domtree.docbook
${DOC}konq-plugins/imgallery.docbook
${DOC}konq-plugins/${C}
${DOC}konq-plugins/${I}
${DOC}konq-plugins/kuick.docbook
${DOC}konq-plugins/mediaplayer.docbook
${DOC}konq-plugins/settings.docbook
${DOC}konq-plugins/uachanger.docbook
${DOC}konq-plugins/validators.docbook
${DOC}konqueror/cmndline.png
${DOC}konqueror/common
${DOC}konqueror/dirtree.png
${DOC}konqueror/dragdrop.png
${DOC}konqueror/filetype1.png
${DOC}konqueror/filetype3.png
${DOC}konqueror/filetype4.png
${DOC}konqueror/${C}
${DOC}konqueror/${I}
${DOC}konqueror/konqorg.png
${DOC}konqueror/parts.png
${DOC}konquest/common
${DOC}konquest/${C}
${DOC}konquest/${I}
${DOC}konsole/common
${DOC}konsole/${C}
${DOC}konsole/${I}
${DOC}konsole/konsole.png
${DOC}kontour/colour.png
${DOC}kontour/common
${DOC}kontour/export.png
${DOC}kontour/${C}
${DOC}kontour/${I}
${DOC}kontour/open_dialog.png
${DOC}kontour/polygon-setup.png
${DOC}kontour/save_dialog.png
${DOC}kooka/common
${DOC}kooka/${C}
${DOC}kooka/${I}
${DOC}korganizer/common
${DOC}korganizer/${C}
${DOC}korganizer/${I}
${DOC}korn/common
${DOC}korn/${C}
${DOC}korn/${I}
${DOC}koshell/common
${DOC}koshell/${C}
${DOC}koshell/${I}
${DOC}kpackage/common
${DOC}kpackage/${C}
${DOC}kpackage/${I}
${DOC}kpager/common
${DOC}kpager/${C}
${DOC}kpager/${I}
${DOC}kpager/screenshot.png
${DOC}kpager/settings.png
${DOC}kpaint/common
${DOC}kpaint/${C}
${DOC}kpaint/${I}
${DOC}kpat/common
${DOC}kpat/${C}
${DOC}kpat/${I}
${DOC}kpat/man.docbook
${DOC}kpf/common
${DOC}kpf/${C}
${DOC}kpf/${I}
${DOC}kpilot/address-app.png
${DOC}kpilot/common
${DOC}kpilot/conduit-knotes.png
${DOC}kpilot/conduit-popmail-kmail.png
${DOC}kpilot/conduit-popmail-recv-method.png
${DOC}kpilot/conduit-popmail-send-as.png
${DOC}kpilot/conduit-popmail-send-method.png
${DOC}kpilot/conduit-popmail-sendmail.png
${DOC}kpilot/conduit-popmail-smtp.png
${DOC}kpilot/conduit-popmail-top.png
${DOC}kpilot/conduit-vcal.png
${DOC}kpilot/file-app.png
${DOC}kpilot/${C}
${DOC}kpilot/${I}
${DOC}kpilot/main-app.png
${DOC}kpilot/memo-app.png
${DOC}kpilot/setup-address.png
${DOC}kpilot/setup-conduit.png
${DOC}kpilot/setup-dbspecial.png
${DOC}kpilot/setup-general.png
${DOC}kpilot/setup-sync.png
${DOC}kpm/common
${DOC}kpm/${C}
${DOC}kpm/${I}
${DOC}kpm/kpmjobs.png
${DOC}kpm/kpmmemory.png
${DOC}kpm/kpmstart.png
${DOC}kpm/kpmtext.png
${DOC}kpoker/common
${DOC}kpoker/${C}
${DOC}kpoker/${I}
${DOC}kpoker/kpoker1.png
${DOC}kpoker/kpoker2.png
${DOC}kppp/accounting.docbook
${DOC}kppp/callback.docbook
${DOC}kppp/chap.docbook
${DOC}kppp/common
${DOC}kppp/dialog-setup.docbook
${DOC}kppp/getting-online.docbook
${DOC}kppp/global-settings.docbook
${DOC}kppp/hayes.docbook
${DOC}kppp/${C}
${DOC}kppp/${I}
${DOC}kppp/kppp-account-accounting-tab.png
${DOC}kppp/kppp-account-dial-tab.png
${DOC}kppp/kppp-account-dns-tab.png
${DOC}kppp/kppp-account-execute-tab.png
${DOC}kppp/kppp-account-gateway-tab.png
${DOC}kppp/kppp-account-ip-tab.png
${DOC}kppp/kppp-account-login-script-tab.png
${DOC}kppp/kppp-config.png
${DOC}kppp/kppp-device-tab.png
${DOC}kppp/kppp-dialler-tab.png
${DOC}kppp/kppp-faq.docbook
${DOC}kppp/kppp-graph-tab.png
${DOC}kppp/kppp-misc-tab.png
${DOC}kppp/kppp-modem-tab.png
${DOC}kppp/kppp-wizard.png
${DOC}kppp/security.docbook
${DOC}kppp/tricks.docbook
${DOC}kppp/wizard.docbook
${DOC}kpresenter/barmenus.png
${DOC}kpresenter/barstyle1.png
${DOC}kpresenter/barstyle2.png
${DOC}kpresenter/barstyle3.png
${DOC}kpresenter/barstyle4.png
${DOC}kpresenter/barstyle5.png
${DOC}kpresenter/barstyle6.png
${DOC}kpresenter/barstyle7.png
${DOC}kpresenter/common
${DOC}kpresenter/faq.docbook
${DOC}kpresenter/great-presentations.docbook
${DOC}kpresenter/guides.docbook
${DOC}kpresenter/htmlshow01.png
${DOC}kpresenter/htmlshow02.png
${DOC}kpresenter/htmlshow03.png
${DOC}kpresenter/htmlshow04.png
${DOC}kpresenter/htmlshow05.png
${DOC}kpresenter/htmlshow07.png
${DOC}kpresenter/${C}
${DOC}kpresenter/${I}
${DOC}kpresenter/menuedit.png
${DOC}kpresenter/menuextra.png
${DOC}kpresenter/menufile.png
${DOC}kpresenter/menuinsert.png
${DOC}kpresenter/menus.docbook
${DOC}kpresenter/menuscreen.png
${DOC}kpresenter/menutext.png
${DOC}kpresenter/menutools.png
${DOC}kpresenter/menuview.png
${DOC}kpresenter/options.docbook
${DOC}kpresenter/screen.docbook
${DOC}kpresenter/settings01.png
${DOC}kpresenter/settings03.png
${DOC}kpresenter/settings04.png
${DOC}kpresenter/settings05.png
${DOC}kpresenter/settings06.png
${DOC}kpresenter/template02.png
${DOC}kpresenter/template03.png
${DOC}kpresenter/template04.png
${DOC}kpresenter/template06.png
${DOC}kpresenter/template07.png
${DOC}kpresenter/textmenu01.png
${DOC}kpresenter/textmenu02.png
${DOC}kpresenter/textmenu03.png
${DOC}kpresenter/textmenu03a.png
${DOC}kpresenter/toolsmenu01.png
${DOC}kpresenter/tut01.png
${DOC}kpresenter/tut02.png
${DOC}kpresenter/tut03.png
${DOC}kpresenter/tut04.png
${DOC}kpresenter/tut05.png
${DOC}kpresenter/tut06.png
${DOC}kpresenter/tut07.png
${DOC}kpresenter/tut08.png
${DOC}kpresenter/tut09.png
${DOC}kpresenter/tut10.png
${DOC}kpresenter/tut11.png
${DOC}kpresenter/tut12.png
${DOC}kpresenter/tut13.png
${DOC}kpresenter/tut14.png
${DOC}kpresenter/tut15.png
${DOC}kpresenter/tut16.png
${DOC}kpresenter/tut17.png
${DOC}kpresenter/tut18.png
${DOC}kpresenter/tut19.png
${DOC}kpresenter/tut20.png
${DOC}kpresenter/tut21.png
${DOC}kpresenter/tut22.png
${DOC}kpresenter/tut23.png
${DOC}kpresenter/tutorial.docbook
${DOC}kreversi/common
${DOC}kreversi/${C}
${DOC}kreversi/${I}
${DOC}kreversi/kreversi1.png
${DOC}kruler/common
${DOC}kruler/${C}
${DOC}kruler/${I}
${DOC}ksame/common
${DOC}ksame/${C}
${DOC}ksame/${I}
${DOC}kscd/common
${DOC}kscd/${C}
${DOC}kscd/${I}
${DOC}kscd/kscd.png
${DOC}kscd/kscd12.png
${DOC}kscd/kscd13.png
${DOC}kscd/kscd14.png
${DOC}kscd/kscd16.png
${DOC}kscd/kscd19.png
${DOC}kscd/kscd2.png
${DOC}kscd/kscd3.png
${DOC}kscore/common
${DOC}kscore/${C}
${DOC}kscore/${I}
${DOC}kshisen/common
${DOC}kshisen/${C}
${DOC}kshisen/${I}
${DOC}ksirc/common
${DOC}ksirc/${C}
${DOC}ksirc/${I}
${DOC}ksirtet/common
${DOC}ksirtet/${C}
${DOC}ksirtet/${I}
${DOC}ksnake/common
${DOC}ksnake/${C}
${DOC}ksnake/${I}
${DOC}ksnapshot/common
${DOC}ksnapshot/${C}
${DOC}ksnapshot/${I}
${DOC}ksnapshot/preview.png
${DOC}ksnapshot/window.png
${DOC}ksokoban/common
${DOC}ksokoban/${C}
${DOC}ksokoban/${I}
${DOC}kspaceduel/common
${DOC}kspaceduel/${C}
${DOC}kspaceduel/${I}
${DOC}kspaceduel/kspaceduel1.png
${DOC}kspaceduel/kspaceduel2.png
${DOC}kspaceduel/kspaceduel3.png
${DOC}kspell/common
${DOC}kspell/${C}
${DOC}kspell/${I}
${DOC}kspread/common
${DOC}kspread/${C}
${DOC}kspread/${I}
${DOC}kstars/ai-contents.docbook
${DOC}kstars/astroinfo.docbook
${DOC}kstars/commands.docbook
${DOC}kstars/common
${DOC}kstars/config.docbook
${DOC}kstars/cpoles.docbook
${DOC}kstars/credits.docbook
${DOC}kstars/csphere.docbook
${DOC}kstars/ecliptic.docbook
${DOC}kstars/equinox.docbook
${DOC}kstars/faq.docbook
${DOC}kstars/geocoords.docbook
${DOC}kstars/greatcircle.docbook
${DOC}kstars/horizon.docbook
${DOC}kstars/hourangle.docbook
${DOC}kstars/${C}
${DOC}kstars/${I}
${DOC}kstars/install.docbook
${DOC}kstars/julianday.docbook
${DOC}kstars/leapyear.docbook
${DOC}kstars/meridian.docbook
${DOC}kstars/precession.docbook
${DOC}kstars/quicktour.docbook
${DOC}kstars/retrograde.docbook
${DOC}kstars/screen1.png
${DOC}kstars/screen2.png
${DOC}kstars/screen3.png
${DOC}kstars/screen4.png
${DOC}kstars/sidereal.docbook
${DOC}kstars/skycoords.docbook
${DOC}kstars/timezones.docbook
${DOC}kstars/utime.docbook
${DOC}kstars/zenith.docbook
${DOC}ksysguard/common
${DOC}ksysguard/${C}
${DOC}ksysguard/${I}
${DOC}ksysv/common
${DOC}ksysv/${C}
${DOC}ksysv/${I}
${DOC}ktalkd/common
${DOC}ktalkd/${C}
${DOC}ktalkd/${I}
${DOC}kteatime/common
${DOC}kteatime/config.png
${DOC}kteatime/${C}
${DOC}kteatime/${I}
${DOC}ktouch/common
${DOC}ktouch/${C}
${DOC}ktouch/${I}
${DOC}ktouch/screenshot1.png
${DOC}ktouch/screenshot2.png
${DOC}ktouch/screenshot3.png
${DOC}ktron/common
${DOC}ktron/${C}
${DOC}ktron/${I}
${DOC}ktuberling/common
${DOC}ktuberling/${C}
${DOC}ktuberling/${I}
${DOC}ktuberling/menu.edit.png
${DOC}ktuberling/menu.file.png
${DOC}ktuberling/menu.help.png
${DOC}ktuberling/menu.option.png
${DOC}ktuberling/menu.raw.png
${DOC}ktuberling/technical-reference.docbook
${DOC}kugar/common
${DOC}kugar/datadtd.docbook
${DOC}kugar/dataref.docbook
${DOC}kugar/${C}
${DOC}kugar/${I}
${DOC}kugar/kugar.png
${DOC}kugar/template-elements.docbook
${DOC}kugar/template.docbook
${DOC}kugar/templatedtd.docbook
${DOC}kuickshow/common
${DOC}kuickshow/${C}
${DOC}kuickshow/${I}
${DOC}kuickshow/screenshot.png
${DOC}kuser/common
${DOC}kuser/${C}
${DOC}kuser/${I}
${DOC}kview/common
${DOC}kview/${C}
${DOC}kview/${I}
${DOC}kview/snapshot1.png
${DOC}kview/snapshot2.png
${DOC}kview/snapshot3.png
${DOC}kview/snapshot4.png
${DOC}kview/snapshot5.png
${DOC}kview/snapshot6.png
${DOC}kview/snapshot7.png
${DOC}kview/snapshot8.png
${DOC}kview/snapshot9.png
${DOC}kvoctrain/art-query-dlg.png
${DOC}kvoctrain/common
${DOC}kvoctrain/comp-query-dlg.png
${DOC}kvoctrain/docprop1-dlg.png
${DOC}kvoctrain/docprop2-dlg.png
${DOC}kvoctrain/docprop6-dlg.png
${DOC}kvoctrain/entry1-dlg.png
${DOC}kvoctrain/entry2-dlg.png
${DOC}kvoctrain/entry3-dlg.png
${DOC}kvoctrain/entry4-dlg.png
${DOC}kvoctrain/entry5-dlg.png
${DOC}kvoctrain/entry6-dlg.png
${DOC}kvoctrain/${C}
${DOC}kvoctrain/${I}
${DOC}kvoctrain/lang1-dlg.png
${DOC}kvoctrain/mainview.png
${DOC}kvoctrain/mu-query-dlg.png
${DOC}kvoctrain/options1-dlg.png
${DOC}kvoctrain/options2-dlg.png
${DOC}kvoctrain/options3-dlg.png
${DOC}kvoctrain/options4-dlg.png
${DOC}kvoctrain/pron-dlg.png
${DOC}kvoctrain/q-opt1-dlg.png
${DOC}kvoctrain/q-opt2-dlg.png
${DOC}kvoctrain/q-opt3-dlg.png
${DOC}kvoctrain/q-opt4-dlg.png
${DOC}kvoctrain/query-dlg.png
${DOC}kvoctrain/stat1-dlg.png
${DOC}kvoctrain/stat2-dlg.png
${DOC}kvoctrain/syn-query-dlg.png
${DOC}kvoctrain/verb-query-dlg.png
${DOC}kweather/common
${DOC}kweather/${C}
${DOC}kweather/${I}
${DOC}kwin4/common
${DOC}kwin4/${C}
${DOC}kwin4/${I}
${DOC}kword/ChooseTempDia.png
${DOC}kword/Tut1.png
${DOC}kword/Tut11a.png
${DOC}kword/Tut11b.png
${DOC}kword/Tut13.png
${DOC}kword/Tut14.png
${DOC}kword/Tut14a.png
${DOC}kword/Tut14b.png
${DOC}kword/Tut15.png
${DOC}kword/Tut15b.png
${DOC}kword/Tut16.png
${DOC}kword/Tut18.png
${DOC}kword/Tut19.png
${DOC}kword/Tut2.png
${DOC}kword/Tut21.png
${DOC}kword/Tut22.png
${DOC}kword/Tut3.png
${DOC}kword/Tut4.png
${DOC}kword/Tut7.png
${DOC}kword/Tut8.png
${DOC}kword/auto1.png
${DOC}kword/auto2.png
${DOC}kword/auto3.png
${DOC}kword/basic.png
${DOC}kword/basics.docbook
${DOC}kword/columns.docbook
${DOC}kword/common
${DOC}kword/ctab2.png
${DOC}kword/delcoldlg.png
${DOC}kword/delrowdlg.png
${DOC}kword/do_not_translate.docbook
${DOC}kword/dtab2.png
${DOC}kword/dtpfmtpg1.png
${DOC}kword/dtpfmtpg2.png
${DOC}kword/editing.docbook
${DOC}kword/fchardlg.png
${DOC}kword/finddlg.png
${DOC}kword/formatchar.docbook
${DOC}kword/formatframes.docbook
${DOC}kword/formatpara.docbook
${DOC}kword/formframe1.png
${DOC}kword/formframe2.png
${DOC}kword/formframe4.png
${DOC}kword/formulas.docbook
${DOC}kword/fpara1.png
${DOC}kword/fpara2.png
${DOC}kword/fpara3.png
${DOC}kword/fpara4.png
${DOC}kword/fpara5.png
${DOC}kword/framers.png
${DOC}kword/frames.docbook
${DOC}kword/fundimentals.docbook
${DOC}kword/graphics.docbook
${DOC}kword/headerfooter.docbook
${DOC}kword/${C}
${DOC}kword/${I}
${DOC}kword/inscoldlg.png
${DOC}kword/insertmisc.docbook
${DOC}kword/insrowdlg.png
${DOC}kword/instab1.png
${DOC}kword/instab2.png
${DOC}kword/intro1.png
${DOC}kword/intro2.png
${DOC}kword/intro3.png
${DOC}kword/kparts.docbook
${DOC}kword/kwordtechinfo.docbook
${DOC}kword/ltab2.png
${DOC}kword/mbtb.docbook
${DOC}kword/obtkb.png
${DOC}kword/obttb.png
${DOC}kword/opendlg.png
${DOC}kword/opt.docbook
${DOC}kword/opt1.png
${DOC}kword/opt2.png
${DOC}kword/optkb.png
${DOC}kword/opttb.png
${DOC}kword/pageformat.docbook
${DOC}kword/pntdlg.png
${DOC}kword/pntdlg1.png
${DOC}kword/repldlg.png
${DOC}kword/rtab2.png
${DOC}kword/ruler.png
${DOC}kword/saved1.png
${DOC}kword/saved2.png
${DOC}kword/savedlg.png
${DOC}kword/savetmpl1.png
${DOC}kword/savetmpl2.png
${DOC}kword/savetmpl3.png
${DOC}kword/savetmpl4.png
${DOC}kword/screen.png
${DOC}kword/select1.png
${DOC}kword/spelldlg.png
${DOC}kword/storeprint.docbook
${DOC}kword/styldlg1.png
${DOC}kword/styldlg2.png
${DOC}kword/styldlg3.png
${DOC}kword/styldlg4.png
${DOC}kword/styldlg5.png
${DOC}kword/styldlg6.png
${DOC}kword/styldlg7.png
${DOC}kword/styldlg8.png
${DOC}kword/styles.docbook
${DOC}kword/table.docbook
${DOC}kword/tabstops.docbook
${DOC}kword/tb2.png
${DOC}kword/tb3.png
${DOC}kword/tb4.png
${DOC}kword/tbmax.png
${DOC}kword/techinfo.docbook
${DOC}kword/templatecreation.docbook
${DOC}kword/toc.docbook
${DOC}kword/tutorial.docbook
${DOC}kword/wpfmtpg1.png
${DOC}kword/wpfmtpg2.png
${DOC}kword/wpfmtpg3.png
${DOC}kworldclock/common
${DOC}kworldclock/${C}
${DOC}kworldclock/${I}
${DOC}kwrite/common
${DOC}kwrite/${C}
${DOC}kwrite/${I}
${DOC}kwuftpd/common
${DOC}kwuftpd/directories.png
${DOC}kwuftpd/${C}
${DOC}kwuftpd/${I}
${DOC}kwuftpd/logging.png
${DOC}kwuftpd/messages.png
${DOC}kwuftpd/ratios.png
${DOC}kwuftpd/security.png
${DOC}kwuftpd/uploads.png
${DOC}kwuftpd/user_classes.png
${DOC}kwuftpd/virtual.png
${DOC}lisa/common
${DOC}lisa/${C}
${DOC}lisa/${I}
${DOC}lskat/common
${DOC}lskat/${C}
${DOC}lskat/${I}
${DOC}noatun/common
${DOC}noatun/${C}
${DOC}noatun/${I}
${DOC}thesaurus/common
${DOC}thesaurus/${C}
${DOC}thesaurus/${I}
${LOC}Kiten.mo
${LOC}aktion.mo
${LOC}amor.mo
${LOC}appletproxy.mo
${LOC}ark.mo
${LOC}artsbuilder.mo
${LOC}artscontrol.mo
${LOC}atlantik.mo
${LOC}atlantikdesigner.mo
${LOC}babelfish.mo
${LOC}caitoo.mo
${LOC}cervisia.mo
${LOC}childpanelextension.mo
${LOC}clockapplet.mo
${LOC}colfind.mo
${LOC}columbo.mo
${LOC}cookbook.mo
${LOC}cupsdconf.mo
${LOC}desktop.mo
${LOC}devcenter.mo
${LOC}dirfilterplugin.mo
${LOC}domtreeviewer.mo
${LOC}drkonqi.mo
${LOC}dub.mo
${LOC}dvd.mo
${LOC}empath.mo
${LOC}extensionproxy.mo
${LOC}filetypes.mo
${LOC}fontinst.mo
${LOC}gideon.mo
${LOC}gofai.mo
${LOC}htmlsearch.mo
${LOC}imagerename_plugin.mo
${LOC}imgalleryplugin.mo
${LOC}kab.mo
${LOC}kab3.mo
${LOC}kaboodle.mo
${LOC}kaccess.mo
${LOC}kaddressbook.mo
${LOC}kafka.mo
${LOC}kalaktic.mo
${LOC}kalarm.mo
${LOC}kalarmd.mo
${LOC}kalarmdgui.mo
${LOC}kandy.mo
${LOC}kaphorism.mo
${LOC}kappfinder.mo
${LOC}karchiver.mo
${LOC}karm.mo
${LOC}kasbarextension.mo
${LOC}kasteroids.mo
${LOC}katalog.mo
${LOC}kate.mo
${LOC}katehelloworld.mo
${LOC}katehtmltools.mo
${LOC}kateinsertcommand.mo
${LOC}kateopenheader.mo
${LOC}katepart.mo
${LOC}kateprojectmanager.mo
${LOC}katetextfilter.mo
${LOC}katexmltools.mo
${LOC}katomic.mo
${LOC}kaudiocreator.mo
${LOC}kautorun.mo
${LOC}kbabel.mo
${LOC}kbackgammon.mo
${LOC}kbattleship.mo
${LOC}kbiff.mo
${LOC}kblackbox.mo
${LOC}kbounce.mo
${LOC}kbugbuster.mo
${LOC}kcalc.mo
${LOC}kcardchooser.mo
${LOC}kcharselect.mo
${LOC}kcharselectapplet.mo
${LOC}kcli.mo
${LOC}kcm_scsimanager.mo
${LOC}kcm_splash.mo
${LOC}kcmaccess.mo
${LOC}kcmarts.mo
${LOC}kcmaudiocd.mo
${LOC}kcmbackground.mo
${LOC}kcmbell.mo
${LOC}kcmbind.mo
${LOC}kcmcddb.mo
${LOC}kcmcolors.mo
${LOC}kcmcrypto.mo
${LOC}kcmcss.mo
${LOC}kcmdhcpd.mo
${LOC}kcmemail.mo
${LOC}kcmenergy.mo
${LOC}kcmfonts.mo
${LOC}kcmgofai.mo
${LOC}kcmhtmlsearch.mo
${LOC}kcmicons.mo
${LOC}kcminfo.mo
${LOC}kcminput.mo
${LOC}kcmioslaveinfo.mo
${LOC}kcmiwatcher.mo
${LOC}kcmkamera.mo
${LOC}kcmkclock.mo
${LOC}kcmkdb.mo
${LOC}kcmkeys.mo
${LOC}kcmkicker.mo
${LOC}kcmkio.mo
${LOC}kcmkmix.mo
${LOC}kcmkonq.mo
${LOC}kcmkonqhtml.mo
${LOC}kcmkonsole.mo
${LOC}kcmktalkd.mo
${LOC}kcmkuick.mo
${LOC}kcmkurifilt.mo
${LOC}kcmkwindecoration.mo
${LOC}kcmkwintheme.mo
${LOC}kcmkwm.mo
${LOC}kcmkxmlrpcd.mo
${LOC}kcmlanbrowser.mo
${LOC}kcmlaptop.mo
${LOC}kcmlaunch.mo
${LOC}kcmlayout.mo
${LOC}kcmlilo.mo
${LOC}kcmlinuz.mo
${LOC}kcmlocale.mo
${LOC}kcmmediacontrol.mo
${LOC}kcmmidi.mo
${LOC}kcmnapster.mo
${LOC}kcmnewsticker.mo
${LOC}kcmnic.mo
${LOC}kcmnotify.mo
${LOC}kcmodbc.mo
${LOC}kcmsamba.mo
${LOC}kcmsblive.mo
${LOC}kcmscreensaver.mo
${LOC}kcmsmartcard.mo
${LOC}kcmsmserver.mo
${LOC}kcmsocks.mo
${LOC}kcmspellchecking.mo
${LOC}kcmstyle.mo
${LOC}kcmtaskbar.mo
${LOC}kcmthemes.mo
${LOC}kcmusb.mo
${LOC}kcmuserenv.mo
${LOC}kcmvdvd.mo
${LOC}kcmwidgetsettings.mo
${LOC}kcoloredit.mo
${LOC}kcontrol.mo
${LOC}kcron.mo
${LOC}kdao.mo
${LOC}kdat.mo
${LOC}kdbbrowser.mo
${LOC}kdcop.mo
${LOC}kdebugdialog.mo
${LOC}kdelibs.mo
${LOC}kdepasswd.mo
${LOC}kdeprintfax.mo
${LOC}kdesktop.mo
${LOC}kdesktop_lock.mo
${LOC}kdessh.mo
${LOC}kdestdifacedemo.mo
${LOC}kdesu.mo
${LOC}kdesud.mo
${LOC}kdevelop.mo
${LOC}kdevtipofday.mo
${LOC}kdf.mo
${LOC}kdict.mo
${LOC}kdictapplet.mo
${LOC}kdmchooser.mo
${LOC}kdmconfig.mo
${LOC}kdmgreet.mo
${LOC}kdvi.mo
${LOC}kedit.mo
${LOC}keduca.mo
${LOC}kenolaba.mo
${LOC}keystone.mo
${LOC}kfax.mo
${LOC}kfifteenapplet.mo
${LOC}kfile_m3u.mo
${LOC}kfile_mp3.mo
${LOC}kfile_ogg.mo
${LOC}kfile_pdf.mo
${LOC}kfile_png.mo
${LOC}kfile_ps.mo
${LOC}kfile_wav.mo
${LOC}kfind.mo
${LOC}kfindpart.mo
${LOC}kfinger.mo
${LOC}kfloppy.mo
${LOC}kfmclient.mo
${LOC}kfmexec.mo
${LOC}kformeditor.mo
${LOC}kformviewer.mo
${LOC}kfortune.mo
${LOC}kfract.mo
${LOC}kgantt.mo
${LOC}kgeo.mo
${LOC}kget.mo
${LOC}kghostview.mo
${LOC}kgnuplot.mo
${LOC}kgrapher.mo
${LOC}khangman.mo
${LOC}khelpcenter.mo
${LOC}khexedit.mo
${LOC}khotkeys.mo
${LOC}khtmlsettingsplugin.mo
${LOC}kicker.mo
${LOC}kiconedit.mo
${LOC}kicq.mo
${LOC}kikbd.mo
${LOC}kim.mo
${LOC}kio_audiocd.mo
${LOC}kio_finger.mo
${LOC}kio_floppy.mo
${LOC}kio_help.mo
${LOC}kio_imap4.mo
${LOC}kio_lan.mo
${LOC}kio_man.mo
${LOC}kio_nfs.mo
${LOC}kio_nntp.mo
${LOC}kio_pop3.mo
${LOC}kio_print.mo
${LOC}kio_sftp.mo
${LOC}kio_smb.mo
${LOC}kio_smbro.mo
${LOC}kio_smtp.mo
${LOC}kit.mo
${LOC}kjobviewer.mo
${LOC}kjots.mo
${LOC}kjumpingcube.mo
${LOC}klaptopdaemon.mo
${LOC}klatin.mo
${LOC}klegacyimport.mo
${LOC}kless.mo
${LOC}klettres.mo
${LOC}klines.mo
${LOC}klipper.mo
${LOC}kljettool.mo
${LOC}klock.mo
${LOC}klpq.mo
${LOC}klprfax.mo
${LOC}kmahjongg.mo
${LOC}kmail.mo
${LOC}kmailcvt.mo
${LOC}kmake.mo
${LOC}kmcop.mo
${LOC}kmenuedit.mo
${LOC}kmessage.mo
${LOC}kmessedwords.mo
${LOC}kmid.mo
${LOC}kmidi.mo
${LOC}kmines.mo
${LOC}kminipagerapplet.mo
${LOC}kmix.mo
${LOC}kmms.mo
${LOC}kmoon.mo
${LOC}knetmgr.mo
${LOC}knewsticker.mo
${LOC}knode.mo
${LOC}knotes.mo
${LOC}knotify.mo
${LOC}knu.mo
${LOC}kodo.mo
${LOC}kolf.mo
${LOC}kolourpicker.mo
${LOC}kompare.mo
${LOC}koncd.mo
${LOC}konqsidebar_mediaplayer.mo
${LOC}konqueror.mo
${LOC}konquest.mo
${LOC}konsole.mo
${LOC}konv.mo
${LOC}kooka.mo
${LOC}kopennap.mo
${LOC}korganizer.mo
${LOC}korn.mo
${LOC}kp.mo
${LOC}kpackage.mo
${LOC}kpager.mo
${LOC}kpaint.mo
${LOC}kpartapp.mo
${LOC}kpartsaver.mo
${LOC}kpat.mo
${LOC}kpercentage.mo
${LOC}kpersonalizer.mo
${LOC}kpf.mo
${LOC}kphone.mo
${LOC}kpilot.mo
${LOC}kpixmap2bitmap.mo
${LOC}kpoker.mo
${LOC}kpovmodeler.mo
${LOC}kpplot.mo
${LOC}kppp.mo
${LOC}kppplogview.mo
${LOC}kprinter.mo
${LOC}kreadconfig.mo
${LOC}kregexpeditor.mo
${LOC}kreversi.mo
${LOC}krn.mo
${LOC}kruler.mo
${LOC}krunapplet.mo
${LOC}ksame.mo
${LOC}kscd.mo
${LOC}kscoreapplet.mo
${LOC}kshisen.mo
${LOC}ksirc.mo
${LOC}ksirtet.mo
${LOC}ksmiletris.mo
${LOC}ksmserver.mo
${LOC}ksnake.mo
${LOC}ksnapshot.mo
${LOC}ksokoban.mo
${LOC}kspaceduel.mo
${LOC}ksplash.mo
${LOC}kstars.mo
${LOC}kstart.mo
${LOC}kstartperf.mo
${LOC}kstockticker.mo
${LOC}ksync.mo
${LOC}ksysctrl.mo
${LOC}ksysguard.mo
${LOC}ksystemtrayapplet.mo
${LOC}ksystraycmd.mo
${LOC}ksystrayproxy.mo
${LOC}ksysv.mo
${LOC}ktables.mo
${LOC}ktalk.mo
${LOC}ktalkd.mo
${LOC}ktaskbarapplet.mo
${LOC}kteatime.mo
${LOC}ktetrinet.mo
${LOC}ktimemon.mo
${LOC}ktimer.mo
${LOC}ktip.mo
${LOC}ktouch.mo
${LOC}ktron.mo
${LOC}ktuberling.mo
${LOC}ktux.mo
${LOC}kue.mo
${LOC}kuick_plugin.mo
${LOC}kuickshow.mo
${LOC}kuser.mo
${LOC}kvalgrind.mo
${LOC}kvidmode.mo
${LOC}kview.mo
${LOC}kviewshell.mo
${LOC}kvoctrain.mo
${LOC}kweather.mo
${LOC}kwin.mo
${LOC}kwin4.mo
${LOC}kwin_b2_config.mo
${LOC}kwin_cde_config.mo
${LOC}kwin_default_config.mo
${LOC}kwin_glow_config.mo
${LOC}kwin_icewm_config.mo
${LOC}kwin_modernsys_config.mo
${LOC}kwin_quartz_config.mo
${LOC}kwintv.mo
${LOC}kwireless.mo
${LOC}kwiz.mo
${LOC}kworldclock.mo
${LOC}kwuftpd.mo
${LOC}kxkb.mo
${LOC}kxmlrpcd.mo
${LOC}kxsconfig.mo
${LOC}libatlantik_network.mo
${LOC}libkcal.mo
${LOC}libkdegames.mo
${LOC}libkdehighscores.mo
${LOC}libkdenetwork.mo
${LOC}libkicker.mo
${LOC}libkickermenu_kdeprint.mo
${LOC}libkonq.mo
${LOC}libkscan.mo
${LOC}libkscreensaver.mo
${LOC}libkwincde_config.mo
${LOC}libkwinglow_config.mo
${LOC}libtaskbar.mo
${LOC}libtaskmanager.mo
${LOC}lockout.mo
${LOC}lskat.mo
${LOC}mediacontrol.mo
${LOC}megami.mo
${LOC}multiplayers.mo
${LOC}naughtyapplet.mo
${LOC}noatun.mo
${LOC}nsplugin.mo
${LOC}passwords.mo
${LOC}ppdtranslations.mo
${LOC}pws.mo
${LOC}quicklauncher.mo
${LOC}secpolicy.mo
${LOC}spy.mo
${LOC}taskbarextension.mo
${LOC}twister.mo
${LOC}uachangerplugin.mo
${LOC}validatorsplugin.mo
${LOC}webarchiver.mo
${LOC}zonedclockapplet.mo
share/locale/sv/charset
share/locale/sv/entry.desktop
share/locale/sv/flag.png
@dirrm share/locale/sv/LC_MESSAGES
@dirrm share/locale/sv
@dirrm ${DOC}thesaurus
@dirrm ${DOC}noatun
@dirrm ${DOC}lskat
@dirrm ${DOC}lisa
@dirrm ${DOC}kwuftpd
@dirrm ${DOC}kwrite
@dirrm ${DOC}kworldclock
@dirrm ${DOC}kword
@dirrm ${DOC}kwin4
@dirrm ${DOC}kweather
@dirrm ${DOC}kvoctrain
@dirrm ${DOC}kview
@dirrm ${DOC}kuser
@dirrm ${DOC}kuickshow
@dirrm ${DOC}kugar
@dirrm ${DOC}ktuberling
@dirrm ${DOC}ktron
@dirrm ${DOC}ktouch
@dirrm ${DOC}kteatime
@dirrm ${DOC}ktalkd
@dirrm ${DOC}ksysv
@dirrm ${DOC}ksysguard
@dirrm ${DOC}kstars
@dirrm ${DOC}kspread
@dirrm ${DOC}kspell
@dirrm ${DOC}kspaceduel
@dirrm ${DOC}ksokoban
@dirrm ${DOC}ksnapshot
@dirrm ${DOC}ksnake
@dirrm ${DOC}ksirtet
@dirrm ${DOC}ksirc
@dirrm ${DOC}kshisen
@dirrm ${DOC}kscore
@dirrm ${DOC}kscd
@dirrm ${DOC}ksame
@dirrm ${DOC}kruler
@dirrm ${DOC}kreversi
@dirrm ${DOC}kpresenter
@dirrm ${DOC}kppp
@dirrm ${DOC}kpoker
@dirrm ${DOC}kpm
@dirrm ${DOC}kpilot
@dirrm ${DOC}kpf
@dirrm ${DOC}kpat
@dirrm ${DOC}kpaint
@dirrm ${DOC}kpager
@dirrm ${DOC}kpackage
@dirrm ${DOC}koshell
@dirrm ${DOC}korn
@dirrm ${DOC}korganizer
@dirrm ${DOC}kooka
@dirrm ${DOC}kontour
@dirrm ${DOC}konsole
@dirrm ${DOC}konquest
@dirrm ${DOC}konqueror
@dirrm ${DOC}konq-plugins
@dirrm ${DOC}koncd
@dirrm ${DOC}koffice
@dirrm ${DOC}kodo
@dirrm ${DOC}knotes
@dirrm ${DOC}knode
@dirrm ${DOC}knewsticker
@dirrm ${DOC}kmoon
@dirrm ${DOC}kmix
@dirrm ${DOC}kmines
@dirrm ${DOC}kmidi
@dirrm ${DOC}kmid
@dirrm ${DOC}kmessedwords
@dirrm ${DOC}kmenuedit
@dirrm ${DOC}kmail
@dirrm ${DOC}klprfax
@dirrm ${DOC}klpq
@dirrm ${DOC}kljettool
@dirrm ${DOC}klipper
@dirrm ${DOC}klines
@dirrm ${DOC}klettres
@dirrm ${DOC}kjumpingcube
@dirrm ${DOC}kjots
@dirrm ${DOC}kit
@dirrm ${DOC}kioslave
@dirrm ${DOC}kiconedit
@dirrm ${DOC}kicker-applets
@dirrm ${DOC}kicker
@dirrm ${DOC}khexedit
@dirrm ${DOC}khelpcenter/visualdict
@dirrm ${DOC}khelpcenter/userguide
@dirrm ${DOC}khelpcenter/quickstart
@dirrm ${DOC}khelpcenter/glossary
@dirrm ${DOC}khelpcenter/faq
@dirrm ${DOC}khelpcenter
@dirrm ${DOC}khangman
@dirrm ${DOC}kghostview
@dirrm ${DOC}kgeo
@dirrm ${DOC}kfract
@dirrm ${DOC}kfouleggs
@dirrm ${DOC}kformula
@dirrm ${DOC}kfloppy
@dirrm ${DOC}kfind
@dirrm ${DOC}kenolaba
@dirrm ${DOC}kedit
@dirrm ${DOC}kdvi
@dirrm ${DOC}kdm
@dirrm ${DOC}kdict
@dirrm ${DOC}kdf
@dirrm ${DOC}kdevelop
@dirrm ${DOC}kdesu
@dirrm ${DOC}kdeprint
@dirrm ${DOC}kdebugdialog
@dirrm ${DOC}kdat
@dirrm ${DOC}kcron
@dirrm ${DOC}kcontrol
@dirrm ${DOC}kcoloredit
@dirrm ${DOC}kcalc
@dirrm ${DOC}kbounce
@dirrm ${DOC}kblackbox
@dirrm ${DOC}kbattleship
@dirrm ${DOC}kbackgammon
@dirrm ${DOC}kbabel
@dirrm ${DOC}katomic
@dirrm ${DOC}kate-plugins
@dirrm ${DOC}kate
@dirrm ${DOC}kasteroids
@dirrm ${DOC}karm
@dirrm ${DOC}kandy
@dirrm ${DOC}kalarm
@dirrm ${DOC}kaddressbook
@dirrm ${DOC}kab
@dirrm ${DOC}common
@dirrm ${DOC}cervisia
@dirrm ${DOC}artsbuilder/images
@dirrm ${DOC}artsbuilder
@dirrm ${DOC}ark
@dirrm ${DOC}amor
@dirrm ${DOC}aktion
@dirrm ${DOC}KRegExpEditor
@dirrm share/doc/HTML/sv
@dirrm share/doc/HTML
@dirrm share/apps/ktuberling/sounds/sv
@dirrm share/apps/ktuberling/sounds
@dirrm share/apps/ktuberling
@dirrm share/apps
