module main

fn main() {
	println('It is not recommended to use "v self" with this packaged version. Please use the source distribution of V if you rely on this functionality')
}
