module main

fn main() {
	println('Use "pkg_add -u v" to update V, or if you want more recent V versions, just from V from source, https://github.com/vlang/v#installing-v-from-source')
	println('If the V package is outdated in OpenBSD -current, please notify the maintainer.')
}
