@comment $OpenBSD: PLIST.sv,v 1.2 2002/12/15 16:21:32 espie Exp $
${DOC}kchart/common
${DOC}kchart/${C}
${DOC}kchart/${I}
${DOC}kformula/additional_fonts1.png
${DOC}kformula/ambiguous-string.png
${DOC}kformula/common
${DOC}kformula/esstix-kfo1.png
${DOC}kformula/esstix-kfo2.png
${DOC}kformula/esstix-kfo3.png
${DOC}kformula/green1.png
${DOC}kformula/green2.png
${DOC}kformula/${C}
${DOC}kformula/${I}
${DOC}kformula/kfontinst-right.png
${DOC}kformula/kfontinst1.png
${DOC}kformula/kfontinst2.png
${DOC}kformula/kfontinst3.png
${DOC}kformula/kfontinst4.png
${DOC}kformula/kfontinst5.png
${DOC}kformula/rk-edit0.png
${DOC}kformula/rk-edit1.png
${DOC}kformula/rk-edit2.png
${DOC}kformula/scilab-edit.png
${DOC}kformula/shortcut0.png
${DOC}kformula/shortcut1.png
${DOC}kformula/toolbars.png
${DOC}koffice/common
${DOC}koffice/${C}
${DOC}koffice/${I}
${DOC}koshell/common
${DOC}koshell/${C}
${DOC}koshell/${I}
${DOC}kpresenter/barmenus.png
${DOC}kpresenter/barstyle1.png
${DOC}kpresenter/barstyle2.png
${DOC}kpresenter/barstyle3.png
${DOC}kpresenter/barstyle4.png
${DOC}kpresenter/barstyle5.png
${DOC}kpresenter/barstyle6.png
${DOC}kpresenter/barstyle7.png
${DOC}kpresenter/common
${DOC}kpresenter/faq.docbook
${DOC}kpresenter/great-presentations.docbook
${DOC}kpresenter/guides.docbook
${DOC}kpresenter/htmlshow01.png
${DOC}kpresenter/htmlshow02.png
${DOC}kpresenter/htmlshow03.png
${DOC}kpresenter/htmlshow04.png
${DOC}kpresenter/htmlshow05.png
${DOC}kpresenter/htmlshow07.png
${DOC}kpresenter/${C}
${DOC}kpresenter/${I}
${DOC}kpresenter/menuedit.png
${DOC}kpresenter/menuextra.png
${DOC}kpresenter/menufile.png
${DOC}kpresenter/menuinsert.png
${DOC}kpresenter/menus.docbook
${DOC}kpresenter/menuscreen.png
${DOC}kpresenter/menutext.png
${DOC}kpresenter/menutools.png
${DOC}kpresenter/menuview.png
${DOC}kpresenter/options.docbook
${DOC}kpresenter/screen.docbook
${DOC}kpresenter/settings01.png
${DOC}kpresenter/settings03.png
${DOC}kpresenter/settings04.png
${DOC}kpresenter/settings05.png
${DOC}kpresenter/settings06.png
${DOC}kpresenter/template02.png
${DOC}kpresenter/template03.png
${DOC}kpresenter/template04.png
${DOC}kpresenter/template06.png
${DOC}kpresenter/template07.png
${DOC}kpresenter/textmenu01.png
${DOC}kpresenter/textmenu02.png
${DOC}kpresenter/textmenu03.png
${DOC}kpresenter/textmenu03a.png
${DOC}kpresenter/toolsmenu01.png
${DOC}kpresenter/tut01.png
${DOC}kpresenter/tut02.png
${DOC}kpresenter/tut03.png
${DOC}kpresenter/tut04.png
${DOC}kpresenter/tut05.png
${DOC}kpresenter/tut06.png
${DOC}kpresenter/tut07.png
${DOC}kpresenter/tut08.png
${DOC}kpresenter/tut09.png
${DOC}kpresenter/tut10.png
${DOC}kpresenter/tut11.png
${DOC}kpresenter/tut12.png
${DOC}kpresenter/tut13.png
${DOC}kpresenter/tut14.png
${DOC}kpresenter/tut15.png
${DOC}kpresenter/tut16.png
${DOC}kpresenter/tut17.png
${DOC}kpresenter/tut18.png
${DOC}kpresenter/tut19.png
${DOC}kpresenter/tut20.png
${DOC}kpresenter/tut21.png
${DOC}kpresenter/tut22.png
${DOC}kpresenter/tut23.png
${DOC}kpresenter/tutorial.docbook
${DOC}kspread/chart1.png
${DOC}kspread/common
${DOC}kspread/copy1.png
${DOC}kspread/${C}
${DOC}kspread/${I}
${DOC}kspread/shortcut1.png
${DOC}kspread/shortcut2.png
${DOC}kspread/sort1.png
${DOC}kspread/starting1.png
${DOC}kugar/add_detail.png
${DOC}kugar/add_detail_footer.png
${DOC}kugar/add_detail_header.png
${DOC}kugar/common
${DOC}kugar/datadtd.docbook
${DOC}kugar/dataref.docbook
${DOC}kugar/designer.docbook
${DOC}kugar/file_new.png
${DOC}kugar/${C}
${DOC}kugar/${I}
${DOC}kugar/kugar.png
${DOC}kugar/progguide.docbook
${DOC}kugar/props.png
${DOC}kugar/starting.docbook
${DOC}kugar/template-elements.docbook
${DOC}kugar/template.docbook
${DOC}kugar/templatedtd.docbook
${DOC}kugar/tut_edit_height.png
${DOC}kugar/tut_empty_report.png
${DOC}kugar/tut_file_new.png
${DOC}kugar/tut_rep_complete.png
${DOC}kugar/tut_rep_generated.png
${DOC}kugar/tut_rep_look1.png
${DOC}kugar/tut_rep_look2.png
${DOC}kugar/tut_set_level.png
${DOC}kugar/tutorial.docbook
${DOC}kword/ChooseTempDia.png
${DOC}kword/Tut1.png
${DOC}kword/Tut11a.png
${DOC}kword/Tut11b.png
${DOC}kword/Tut13.png
${DOC}kword/Tut14.png
${DOC}kword/Tut14a.png
${DOC}kword/Tut14b.png
${DOC}kword/Tut15.png
${DOC}kword/Tut15b.png
${DOC}kword/Tut16.png
${DOC}kword/Tut18.png
${DOC}kword/Tut19.png
${DOC}kword/Tut2.png
${DOC}kword/Tut21.png
${DOC}kword/Tut22.png
${DOC}kword/Tut3.png
${DOC}kword/Tut4.png
${DOC}kword/Tut7.png
${DOC}kword/Tut8.png
${DOC}kword/auto1.png
${DOC}kword/auto2.png
${DOC}kword/auto3.png
${DOC}kword/auto4.png
${DOC}kword/autocompdlg.png
${DOC}kword/basic.png
${DOC}kword/basics.docbook
${DOC}kword/bookmarks.docbook
${DOC}kword/bordtb.png
${DOC}kword/colorseldlg.png
${DOC}kword/columns.docbook
${DOC}kword/common
${DOC}kword/ctab2.png
${DOC}kword/delcoldlg.png
${DOC}kword/delrowdlg.png
${DOC}kword/do_not_translate.docbook
${DOC}kword/doccomments.docbook
${DOC}kword/doclinks.docbook
${DOC}kword/docstruct.docbook
${DOC}kword/docstruct.png
${DOC}kword/docvariables.docbook
${DOC}kword/dtab2.png
${DOC}kword/dtpfmtpg1.png
${DOC}kword/dtpfmtpg2.png
${DOC}kword/editing.docbook
${DOC}kword/expression.png
${DOC}kword/expressions.docbook
${DOC}kword/exst.png
${DOC}kword/exul.png
${DOC}kword/fchardlg.png
${DOC}kword/fchardlg2.png
${DOC}kword/finddlg.png
${DOC}kword/finddlg2.png
${DOC}kword/footcfg1.png
${DOC}kword/footcfg3.png
${DOC}kword/footendnotes.docbook
${DOC}kword/formatchar.docbook
${DOC}kword/formatframes.docbook
${DOC}kword/formatpara.docbook
${DOC}kword/formframe1.png
${DOC}kword/formframe2.png
${DOC}kword/formframe3.png
${DOC}kword/formframe4.png
${DOC}kword/formframe5.png
${DOC}kword/formulas.docbook
${DOC}kword/fpara1.png
${DOC}kword/fpara2.png
${DOC}kword/fpara3.png
${DOC}kword/fpara4.png
${DOC}kword/fpara5.png
${DOC}kword/fpara6.png
${DOC}kword/framers.png
${DOC}kword/frames.docbook
${DOC}kword/framestylist.png
${DOC}kword/fundimentals.docbook
${DOC}kword/graphics.docbook
${DOC}kword/headerfooter.docbook
${DOC}kword/${C}
${DOC}kword/${I}
${DOC}kword/inscoldlg.png
${DOC}kword/insdate.png
${DOC}kword/insertfile.docbook
${DOC}kword/insertmisc.docbook
${DOC}kword/insgrph1.png
${DOC}kword/insgrph2.png
${DOC}kword/insrowdlg.png
${DOC}kword/instab1.png
${DOC}kword/instab2.png
${DOC}kword/instime.png
${DOC}kword/intro1.png
${DOC}kword/intro2.png
${DOC}kword/intro3.png
${DOC}kword/kparts.docbook
${DOC}kword/linkdlg.png
${DOC}kword/listdepth1.png
${DOC}kword/listdepth2.png
${DOC}kword/listdepth3.png
${DOC}kword/lists.docbook
${DOC}kword/ltab2.png
${DOC}kword/mailmerge.docbook
${DOC}kword/mbtb.docbook
${DOC}kword/mmerge1.png
${DOC}kword/mmerge2.png
${DOC}kword/mmergesql1.png
${DOC}kword/mmergesql2.png
${DOC}kword/obtkb.png
${DOC}kword/obttb.png
${DOC}kword/opendlg.png
${DOC}kword/opt.docbook
${DOC}kword/opt1.png
${DOC}kword/opt2.png
${DOC}kword/opt3.png
${DOC}kword/opt4.png
${DOC}kword/opt5.png
${DOC}kword/optkb.png
${DOC}kword/optkb2.png
${DOC}kword/opttb.png
${DOC}kword/pageformat.docbook
${DOC}kword/pntdlg.png
${DOC}kword/pntdlg1.png
${DOC}kword/repldlg.png
${DOC}kword/rtab2.png
${DOC}kword/ruler.png
${DOC}kword/saved1.png
${DOC}kword/saved2.png
${DOC}kword/savedlg.png
${DOC}kword/savetmpl1.png
${DOC}kword/savetmpl2.png
${DOC}kword/savetmpl3.png
${DOC}kword/savetmpl4.png
${DOC}kword/screen.png
${DOC}kword/select1.png
${DOC}kword/spelldlg.png
${DOC}kword/storeprint.docbook
${DOC}kword/styldlg1.png
${DOC}kword/styldlg2.png
${DOC}kword/styldlg3.png
${DOC}kword/styldlg4.png
${DOC}kword/styldlg5.png
${DOC}kword/styldlg6.png
${DOC}kword/styldlg7.png
${DOC}kword/styldlg8.png
${DOC}kword/styles.docbook
${DOC}kword/table.docbook
${DOC}kword/tableprop1.png
${DOC}kword/tableprop2.png
${DOC}kword/tablestylist.png
${DOC}kword/tabstops.docbook
${DOC}kword/tb2.png
${DOC}kword/tb3.png
${DOC}kword/tb4.png
${DOC}kword/tblsty.png
${DOC}kword/tbmax.png
${DOC}kword/techinfo.docbook
${DOC}kword/tedittb.png
${DOC}kword/templatecreation.docbook
${DOC}kword/textstyex.png
${DOC}kword/thesaurus.png
${DOC}kword/toc.docbook
${DOC}kword/tutorial.docbook
${DOC}kword/wpfmtpg1.png
${DOC}kword/wpfmtpg2.png
${DOC}kword/wpfmtpg3.png
${DOC}thesaurus/common
${DOC}thesaurus/${C}
${DOC}thesaurus/${I}
${LOC}csvfilter.mo
${LOC}desktop_koffice.mo
${LOC}example.mo
${LOC}graphite.mo
${LOC}karbon.mo
${LOC}kchart.mo
${LOC}kfile_koffice.mo
${LOC}kformula.mo
${LOC}kformulalatexfilter.mo
${LOC}kformulapngfilter.mo
${LOC}kivio.mo
${LOC}koconverter.mo
${LOC}kocryptfilter.mo
${LOC}koffice.mo
${LOC}kontour.mo
${LOC}koshell.mo
${LOC}kounavail.mo
${LOC}kplato.mo
${LOC}kpresenter.mo
${LOC}kpresenterkwordfilter.mo
${LOC}krita.mo
${LOC}kscan_plugin.mo
${LOC}kspread.mo
${LOC}kspreadcalc_calc.mo
${LOC}kspreadqprofilter.mo
${LOC}kthesaurus.mo
${LOC}kugar.mo
${LOC}kword.mo
${LOC}kwordasciifilter.mo
${LOC}kwordhtmlexportfilter.mo
${LOC}kwordhtmlimportfilter.mo
${LOC}kwordlatexfilter.mo
${LOC}kwordmswritefilter.mo
${LOC}olefilterswinword97filter.mo
${LOC}thesaurus_tool.mo
${LOC}xsltexportfilter.mo
${LOC}xsltimportfilter.mo
@dirrm share/locale/sv/LC_MESSAGES
@dirrm share/locale/sv
@dirrm share/locale
@dirrm ${DOC}thesaurus
@dirrm ${DOC}kword
@dirrm ${DOC}kugar
@dirrm ${DOC}kspread
@dirrm ${DOC}kpresenter
@dirrm ${DOC}koshell
@dirrm ${DOC}koffice
@dirrm ${DOC}kformula
@dirrm ${DOC}kchart
@dirrm share/doc/HTML/sv
@dirrm share/doc/HTML
