@comment $OpenBSD: PLIST.sv,v 1.14 2004/02/07 12:29:13 espie Exp $
share/apps/ktuberling/sounds/sv/brosch.wav
share/apps/ktuberling/sounds/sv/cigarr.wav
share/apps/ktuberling/sounds/sv/fluga.wav
share/apps/ktuberling/sounds/sv/glasogon.wav
share/apps/ktuberling/sounds/sv/halsband.wav
share/apps/ktuberling/sounds/sv/halsduk.wav
share/apps/ktuberling/sounds/sv/har.wav
share/apps/ktuberling/sounds/sv/hatt.wav
share/apps/ktuberling/sounds/sv/horn.wav
share/apps/ktuberling/sounds/sv/klocka.wav
share/apps/ktuberling/sounds/sv/mun.wav
share/apps/ktuberling/sounds/sv/mustasch.wav
share/apps/ktuberling/sounds/sv/nasa.wav
share/apps/ktuberling/sounds/sv/oga.wav
share/apps/ktuberling/sounds/sv/ogonbryn.wav
share/apps/ktuberling/sounds/sv/ora.wav
share/apps/ktuberling/sounds/sv/orhange.wav
share/apps/ktuberling/sounds/sv/pingvin.wav
share/apps/ktuberling/sounds/sv/potatismannen.wav
share/apps/ktuberling/sounds/sv/rosett.wav
share/apps/ktuberling/sounds/sv/slips.wav
share/apps/ktuberling/sounds/sv/solglasogon.wav
${DOC}KRegExpEditor/altntool.png
${DOC}KRegExpEditor/anychartool.png
${DOC}KRegExpEditor/boundarytools.png
${DOC}KRegExpEditor/charactertool.png
${DOC}KRegExpEditor/common
${DOC}KRegExpEditor/compoundtool.png
${DOC}KRegExpEditor/${C}
${DOC}KRegExpEditor/${I}
${DOC}KRegExpEditor/linestartendtool.png
${DOC}KRegExpEditor/lookaheadtools.png
${DOC}KRegExpEditor/repeattool.png
${DOC}KRegExpEditor/theEditor.png
${DOC}amor/common
${DOC}amor/${C}
${DOC}amor/${I}
${DOC}ark/common
${DOC}ark/${C}
${DOC}ark/${I}
${DOC}artsbuilder/apis.docbook
${DOC}artsbuilder/arts-structure.png
${DOC}artsbuilder/artsbuilder.docbook
${DOC}artsbuilder/common
${DOC}artsbuilder/detail.docbook
${DOC}artsbuilder/digitalaudio.docbook
${DOC}artsbuilder/faq.docbook
${DOC}artsbuilder/future.docbook
${DOC}artsbuilder/glossary.docbook
${DOC}artsbuilder/gui.docbook
${DOC}artsbuilder/helping.docbook
${DOC}artsbuilder/images/Synth_AMAN_PLAY.png
${DOC}artsbuilder/images/Synth_AMAN_RECORD.png
${DOC}artsbuilder/images/Synth_BRICKWALL_LIMITER.png
${DOC}artsbuilder/images/Synth_CAPTURE.png
${DOC}artsbuilder/images/Synth_DATA.png
${DOC}artsbuilder/images/Synth_FREEVERB.png
${DOC}artsbuilder/images/Synth_FX_CFLANGER.png
${DOC}artsbuilder/images/Synth_MIDI_TEST.png
${DOC}artsbuilder/images/Synth_MOOG_VCF.png
${DOC}artsbuilder/images/Synth_MULTI_ADD.png
${DOC}artsbuilder/images/Synth_NOISE.png
${DOC}artsbuilder/images/Synth_PITCH_SHIFT.png
${DOC}artsbuilder/images/Synth_RECORD.png
${DOC}artsbuilder/images/Synth_TREMOLO.png
${DOC}artsbuilder/images/Synth_WAVE_PULSE.png
${DOC}artsbuilder/images/Synth_WAVE_SOFTSAW.png
${DOC}artsbuilder/${C}
${DOC}artsbuilder/${I}
${DOC}artsbuilder/mcop.docbook
${DOC}artsbuilder/midi.docbook
${DOC}artsbuilder/midiintro.docbook
${DOC}artsbuilder/modules.docbook
${DOC}artsbuilder/porting.docbook
${DOC}artsbuilder/references.docbook
${DOC}artsbuilder/tools.docbook
${DOC}atlantik/common
${DOC}atlantik/${C}
${DOC}atlantik/${I}
${DOC}cervisia/checkout.png
${DOC}cervisia/commit.png
${DOC}cervisia/common
${DOC}cervisia/diff.png
${DOC}cervisia/history.png
${DOC}cervisia/import.png
${DOC}cervisia/${C}
${DOC}cervisia/${I}
${DOC}cervisia/logtree.png
${DOC}cervisia/mainview.png
${DOC}cervisia/resolve.png
${DOC}cervisia/updatetag.png
${DOC}common/1.png
${DOC}common/10.png
${DOC}common/2.png
${DOC}common/3.png
${DOC}common/4.png
${DOC}common/5.png
${DOC}common/6.png
${DOC}common/7.png
${DOC}common/8.png
${DOC}common/9.png
${DOC}common/appheader.html
${DOC}common/artistic-license.html
${DOC}common/bottom1.png
${DOC}common/bottom2.png
${DOC}common/bsd-license.html
${DOC}common/docheadergears.png
${DOC}common/doctop1.png
${DOC}common/doctop1a.png
${DOC}common/doctop1b.png
${DOC}common/doctop2.png
${DOC}common/doxygen.css
${DOC}common/fdl-license
${DOC}common/fdl-license.html
${DOC}common/fdl-translated.html
${DOC}common/footer.html
${DOC}common/gpl-license
${DOC}common/gpl-license.html
${DOC}common/gpl-translated.html
${DOC}common/grad.png
${DOC}common/header.html
${DOC}common/headerbg.png
${DOC}common/kde-common.css
${DOC}common/kde-default.css
${DOC}common/kde-localised.css
${DOC}common/kde-localised.css.template
${DOC}common/kde-web.css
${DOC}common/kde_logo.png
${DOC}common/kde_logo_bg.png
${DOC}common/kmenu.png
${DOC}common/lgpl-license
${DOC}common/lgpl-license.html
${DOC}common/lgpl-translated.html
${DOC}common/logotp3.png
${DOC}common/mainfooter.html
${DOC}common/mainheader.html
${DOC}common/qpl-license.html
${DOC}common/shadow.png
${DOC}common/web-docbottom.png
${DOC}common/web-doctop.png
${DOC}common/x11-license.html
${DOC}common/xml.dcl
${DOC}flashkard/common
${DOC}flashkard/flashkard1.png
${DOC}flashkard/flashkard2.png
${DOC}flashkard/flashkard3.png
${DOC}flashkard/flashkard4.png
${DOC}flashkard/${C}
${DOC}flashkard/${I}
${DOC}juk/common
${DOC}juk/${C}
${DOC}juk/${I}
${DOC}kaboodle/common
${DOC}kaboodle/${C}
${DOC}kaboodle/${I}
${DOC}kaddressbook/common
${DOC}kaddressbook/conf.png
${DOC}kaddressbook/contactdlg.png
${DOC}kaddressbook/exportdlg.png
${DOC}kaddressbook/extension.png
${DOC}kaddressbook/filtereditdlg.png
${DOC}kaddressbook/${C}
${DOC}kaddressbook/${I}
${DOC}kaddressbook/mainwin.png
${DOC}kaddressbook/resourcedlg.png
${DOC}kaddressbook/vieweditdlg.png
${DOC}kalarm/alarmmessage.png
${DOC}kalarm/common
${DOC}kalarm/editwindow.png
${DOC}kalarm/${C}
${DOC}kalarm/${I}
${DOC}kalarm/mainwindow.png
${DOC}kalzium/common
${DOC}kalzium/${C}
${DOC}kalzium/${I}
${DOC}kalzium/screenshot1.png
${DOC}kalzium/screenshot2.png
${DOC}kalzium/screenshot3.png
${DOC}kalzium/settings.png
${DOC}kamera/common
${DOC}kamera/${C}
${DOC}kamera/${I}
${DOC}kandy/common
${DOC}kandy/${C}
${DOC}kandy/${I}
${DOC}karm/common
${DOC}karm/${C}
${DOC}karm/${I}
${DOC}kasteroids/common
${DOC}kasteroids/${C}
${DOC}kasteroids/${I}
${DOC}kate-plugins/common
${DOC}kate-plugins/htmltools.docbook
${DOC}kate-plugins/${C}
${DOC}kate-plugins/${I}
${DOC}kate-plugins/insertcommand.docbook
${DOC}kate-plugins/openheader.docbook
${DOC}kate-plugins/projectmanager.docbook
${DOC}kate-plugins/textfilter.docbook
${DOC}kate-plugins/xmlcheck.docbook
${DOC}kate-plugins/xmltools.docbook
${DOC}kate/advanced.docbook
${DOC}kate/common
${DOC}kate/configdialog01.png
${DOC}kate/configdialog02.png
${DOC}kate/configuring.docbook
${DOC}kate/fundamentals.docbook
${DOC}kate/highlighting.docbook
${DOC}kate/${C}
${DOC}kate/${I}
${DOC}kate/kate.png
${DOC}kate/mdi.docbook
${DOC}kate/menus.docbook
${DOC}kate/mimetypechooser.png
${DOC}kate/part.docbook
${DOC}kate/plugins.docbook
${DOC}kate/regular-expressions.docbook
${DOC}katomic/common
${DOC}katomic/${C}
${DOC}katomic/${I}
${DOC}kbabel/catman.docbook
${DOC}kbabel/common
${DOC}kbabel/dbcan.png
${DOC}kbabel/dictionaries.docbook
${DOC}kbabel/faq.docbook
${DOC}kbabel/glossary.docbook
${DOC}kbabel/${C}
${DOC}kbabel/${I}
${DOC}kbabel/kbabeldict.docbook
${DOC}kbabel/menu.docbook
${DOC}kbabel/preferences.docbook
${DOC}kbabel/roughtranslation.png
${DOC}kbabel/snap1.png
${DOC}kbabel/snap_catalogmanager.png
${DOC}kbabel/snap_kbabeldict.png
${DOC}kbabel/snap_kbabeldict2.png
${DOC}kbabel/using.docbook
${DOC}kbackgammon/common
${DOC}kbackgammon/${C}
${DOC}kbackgammon/${I}
${DOC}kbattleship/common
${DOC}kbattleship/${C}
${DOC}kbattleship/${I}
${DOC}kblackbox/common
${DOC}kblackbox/${C}
${DOC}kblackbox/${I}
${DOC}kbounce/common
${DOC}kbounce/${C}
${DOC}kbounce/${I}
${DOC}kbounce/jezball_corridor1.png
${DOC}kbounce/jezball_corridor2.png
${DOC}kbounce/jezball_newWall.png
${DOC}kbruch/checked.png
${DOC}kbruch/common
${DOC}kbruch/gui_main.png
${DOC}kbruch/${C}
${DOC}kbruch/${I}
${DOC}kbruch/reduced.png
${DOC}kbugbuster/common
${DOC}kbugbuster/${C}
${DOC}kbugbuster/${I}
${DOC}kcachegrind/common
${DOC}kcachegrind/${C}
${DOC}kcachegrind/${I}
${DOC}kcalc/common
${DOC}kcalc/${C}
${DOC}kcalc/${I}
${DOC}kcharselect/common
${DOC}kcharselect/${C}
${DOC}kcharselect/${I}
${DOC}kcoloredit/common
${DOC}kcoloredit/${C}
${DOC}kcoloredit/${I}
${DOC}kcontrol/arts/common
${DOC}kcontrol/arts/${C}
${DOC}kcontrol/arts/${I}
${DOC}kcontrol/arts/midi.docbook
${DOC}kcontrol/background/common
${DOC}kcontrol/background/${C}
${DOC}kcontrol/background/${I}
${DOC}kcontrol/bell/common
${DOC}kcontrol/bell/${C}
${DOC}kcontrol/bell/${I}
${DOC}kcontrol/cache/common
${DOC}kcontrol/cache/${C}
${DOC}kcontrol/cache/${I}
${DOC}kcontrol/clock/common
${DOC}kcontrol/clock/${C}
${DOC}kcontrol/clock/${I}
${DOC}kcontrol/colors/common
${DOC}kcontrol/colors/${C}
${DOC}kcontrol/colors/${I}
${DOC}kcontrol/common
${DOC}kcontrol/cookies/common
${DOC}kcontrol/cookies/${C}
${DOC}kcontrol/cookies/${I}
${DOC}kcontrol/crypto/common
${DOC}kcontrol/crypto/${C}
${DOC}kcontrol/crypto/${I}
${DOC}kcontrol/desktop/common
${DOC}kcontrol/desktop/${C}
${DOC}kcontrol/desktop/${I}
${DOC}kcontrol/desktopbehavior/common
${DOC}kcontrol/desktopbehavior/${C}
${DOC}kcontrol/desktopbehavior/${I}
${DOC}kcontrol/ebrowsing/common
${DOC}kcontrol/ebrowsing/${C}
${DOC}kcontrol/ebrowsing/${I}
${DOC}kcontrol/email/common
${DOC}kcontrol/email/${C}
${DOC}kcontrol/email/${I}
${DOC}kcontrol/energy/common
${DOC}kcontrol/energy/${C}
${DOC}kcontrol/energy/${I}
${DOC}kcontrol/filemanager/common
${DOC}kcontrol/filemanager/${C}
${DOC}kcontrol/filemanager/${I}
${DOC}kcontrol/filemanager/kfileman1.png
${DOC}kcontrol/filemanager/kfileman2.png
${DOC}kcontrol/filetypes/common
${DOC}kcontrol/filetypes/${C}
${DOC}kcontrol/filetypes/${I}
${DOC}kcontrol/fonts/common
${DOC}kcontrol/fonts/${C}
${DOC}kcontrol/fonts/${I}
${DOC}kcontrol/helpindex/common
${DOC}kcontrol/helpindex/${C}
${DOC}kcontrol/helpindex/${I}
${DOC}kcontrol/icons/common
${DOC}kcontrol/icons/${C}
${DOC}kcontrol/icons/${I}
${DOC}kcontrol/${C}
${DOC}kcontrol/${I}
${DOC}kcontrol/kalarmd/common
${DOC}kcontrol/kalarmd/${C}
${DOC}kcontrol/kalarmd/${I}
${DOC}kcontrol/kcmaccess/common
${DOC}kcontrol/kcmaccess/${C}
${DOC}kcontrol/kcmaccess/${I}
${DOC}kcontrol/kcmcss/common
${DOC}kcontrol/kcmcss/${C}
${DOC}kcontrol/kcmcss/${I}
${DOC}kcontrol/kcmfontinst/common
${DOC}kcontrol/kcmfontinst/${C}
${DOC}kcontrol/kcmfontinst/${I}
${DOC}kcontrol/kcmkonsole/common
${DOC}kcontrol/kcmkonsole/${C}
${DOC}kcontrol/kcmkonsole/${I}
${DOC}kcontrol/kcmktalkd/common
${DOC}kcontrol/kcmktalkd/${C}
${DOC}kcontrol/kcmktalkd/${I}
${DOC}kcontrol/kcmlaunch/common
${DOC}kcontrol/kcmlaunch/${C}
${DOC}kcontrol/kcmlaunch/${I}
${DOC}kcontrol/kcmlowbatcrit/common
${DOC}kcontrol/kcmlowbatcrit/${C}
${DOC}kcontrol/kcmlowbatcrit/${I}
${DOC}kcontrol/kcmlowbatwarn/common
${DOC}kcontrol/kcmlowbatwarn/${C}
${DOC}kcontrol/kcmlowbatwarn/${I}
${DOC}kcontrol/kcmnotify/common
${DOC}kcontrol/kcmnotify/${C}
${DOC}kcontrol/kcmnotify/${I}
${DOC}kcontrol/kcmsmserver/common
${DOC}kcontrol/kcmsmserver/${C}
${DOC}kcontrol/kcmsmserver/${I}
${DOC}kcontrol/kcmstyle/common
${DOC}kcontrol/kcmstyle/${C}
${DOC}kcontrol/kcmstyle/${I}
${DOC}kcontrol/kcmtaskbar/common
${DOC}kcontrol/kcmtaskbar/${C}
${DOC}kcontrol/kcmtaskbar/${I}
${DOC}kcontrol/kdm/common
${DOC}kcontrol/kdm/${C}
${DOC}kcontrol/kdm/${I}
${DOC}kcontrol/keyboard/common
${DOC}kcontrol/keyboard/${C}
${DOC}kcontrol/keyboard/${I}
${DOC}kcontrol/keys/common
${DOC}kcontrol/keys/${C}
${DOC}kcontrol/keys/${I}
${DOC}kcontrol/khtml/common
${DOC}kcontrol/khtml/${C}
${DOC}kcontrol/khtml/${I}
${DOC}kcontrol/khtml/nsplugin.docbook
${DOC}kcontrol/kmixcfg/common
${DOC}kcontrol/kmixcfg/${C}
${DOC}kcontrol/kmixcfg/${I}
${DOC}kcontrol/kthememgr/common
${DOC}kcontrol/kthememgr/${C}
${DOC}kcontrol/kthememgr/${I}
${DOC}kcontrol/kwindecoration/common
${DOC}kcontrol/kwindecoration/${C}
${DOC}kcontrol/kwindecoration/${I}
${DOC}kcontrol/kxmlrpcd/common
${DOC}kcontrol/kxmlrpcd/${C}
${DOC}kcontrol/kxmlrpcd/${I}
${DOC}kcontrol/lanbrowser/common
${DOC}kcontrol/lanbrowser/${C}
${DOC}kcontrol/lanbrowser/${I}
${DOC}kcontrol/language/common
${DOC}kcontrol/language/${C}
${DOC}kcontrol/language/${I}
${DOC}kcontrol/laptop/common
${DOC}kcontrol/laptop/${C}
${DOC}kcontrol/laptop/${I}
${DOC}kcontrol/mouse/common
${DOC}kcontrol/mouse/${C}
${DOC}kcontrol/mouse/${I}
${DOC}kcontrol/netpref/common
${DOC}kcontrol/netpref/${C}
${DOC}kcontrol/netpref/${I}
${DOC}kcontrol/panel/common
${DOC}kcontrol/panel/${C}
${DOC}kcontrol/panel/${I}
${DOC}kcontrol/panelappearance/common
${DOC}kcontrol/panelappearance/${C}
${DOC}kcontrol/panelappearance/${I}
${DOC}kcontrol/passwords/common
${DOC}kcontrol/passwords/${C}
${DOC}kcontrol/passwords/${I}
${DOC}kcontrol/powerctrl/common
${DOC}kcontrol/powerctrl/${C}
${DOC}kcontrol/powerctrl/${I}
${DOC}kcontrol/proxy/common
${DOC}kcontrol/proxy/${C}
${DOC}kcontrol/proxy/${I}
${DOC}kcontrol/proxy/socks.docbook
${DOC}kcontrol/screensaver/common
${DOC}kcontrol/screensaver/${C}
${DOC}kcontrol/screensaver/${I}
${DOC}kcontrol/screenshot.png
${DOC}kcontrol/smb/common
${DOC}kcontrol/smb/${C}
${DOC}kcontrol/smb/${I}
${DOC}kcontrol/spellchecking/common
${DOC}kcontrol/spellchecking/${C}
${DOC}kcontrol/spellchecking/${I}
${DOC}kcontrol/useragent/common
${DOC}kcontrol/useragent/${C}
${DOC}kcontrol/useragent/${I}
${DOC}kcontrol/windowmanagement/common
${DOC}kcontrol/windowmanagement/${C}
${DOC}kcontrol/windowmanagement/${I}
${DOC}kcron/common
${DOC}kcron/${C}
${DOC}kcron/${I}
${DOC}kcron/kcron.png
${DOC}kcron/kcronstart.png
${DOC}kcron/newtask.png
${DOC}kcron/newvariable.png
${DOC}kcron/print.png
${DOC}kdat/common
${DOC}kdat/${C}
${DOC}kdat/${I}
${DOC}kdebugdialog/common
${DOC}kdebugdialog/${C}
${DOC}kdebugdialog/${I}
${DOC}kdeprint/add-printer-wiz.docbook
${DOC}kdeprint/common
${DOC}kdeprint/cups-config.docbook
${DOC}kdeprint/cups-filterarchitecture-kivio-70Percent-scaled.png
${DOC}kdeprint/cupsaddprinterwizard1.png
${DOC}kdeprint/cupsaddprinterwizard2_backendselection.png
${DOC}kdeprint/cupsaddprinterwizard3_networkscan.png
${DOC}kdeprint/cupsaddprinterwizard4_networkscan_config.png
${DOC}kdeprint/cupsoptions.docbook
${DOC}kdeprint/cupsserverconfiguration1_welcome.png
${DOC}kdeprint/extensions.docbook
${DOC}kdeprint/external-command.docbook
${DOC}kdeprint/final-word.docbook
${DOC}kdeprint/getting-started.docbook
${DOC}kdeprint/highlights.docbook
${DOC}kdeprint/${C}
${DOC}kdeprint/${I}
${DOC}kdeprint/kcontrolcenter-printmanager-jobcontrol-2.png
${DOC}kdeprint/kcron_to_be_printed.png
${DOC}kdeprint/kdeprint-jobviewer.png
${DOC}kdeprint/kprinter-as-netscape-printcommand.png
${DOC}kdeprint/kprinter-kivio.png
${DOC}kdeprint/kprinter.png
${DOC}kdeprint/kprinter_called_from_run_command.png
${DOC}kdeprint/kprinter_with_kcron_developer_special.png
${DOC}kdeprint/lpd.docbook
${DOC}kdeprint/lpr-bsd.docbook
${DOC}kdeprint/lprng.docbook
${DOC}kdeprint/rlpr.docbook
${DOC}kdeprint/steinbruch_scaled.png
${DOC}kdeprint/tech-overview.docbook
${DOC}kdeprint/theory.docbook
${DOC}kdesu/common
${DOC}kdesu/${C}
${DOC}kdesu/${I}
${DOC}kdf/common
${DOC}kdf/${C}
${DOC}kdf/${I}
${DOC}kdf/kdf.png
${DOC}kdf/kdf_config.png
${DOC}kdict/applet.png
${DOC}kdict/common
${DOC}kdict/conf.png
${DOC}kdict/${C}
${DOC}kdict/${I}
${DOC}kdict/mainwin.png
${DOC}kdict/seteditor.png
${DOC}kdm/common
${DOC}kdm/${C}
${DOC}kdm/${I}
${DOC}kdm/kdmrc-ref.docbook
${DOC}kdvi/common
${DOC}kdvi/${C}
${DOC}kdvi/${I}
${DOC}kdvi/optionrequester1.png
${DOC}kdvi/optionrequester2.png
${DOC}kedit/common
${DOC}kedit/${C}
${DOC}kedit/${I}
${DOC}keduca/common
${DOC}keduca/${C}
${DOC}keduca/${I}
${DOC}keduca/screenshot.png
${DOC}kenolaba/common
${DOC}kenolaba/${C}
${DOC}kenolaba/${I}
${DOC}kfind/common
${DOC}kfind/${C}
${DOC}kfind/${I}
${DOC}kfloppy/common
${DOC}kfloppy/${C}
${DOC}kfloppy/${I}
${DOC}kfouleggs/common
${DOC}kfouleggs/gamescreen.png
${DOC}kfouleggs/${C}
${DOC}kfouleggs/${I}
${DOC}kgamma/common
${DOC}kgamma/${C}
${DOC}kgamma/${I}
${DOC}kget/common
${DOC}kget/cr22-action-tool_delay.png
${DOC}kget/cr22-action-tool_disconnect.png
${DOC}kget/cr22-action-tool_drop_target.png
${DOC}kget/cr22-action-tool_expert.png
${DOC}kget/cr22-action-tool_logwindow.png
${DOC}kget/cr22-action-tool_offline_mode_off.png
${DOC}kget/cr22-action-tool_offline_mode_on.png
${DOC}kget/cr22-action-tool_paste.png
${DOC}kget/cr22-action-tool_pause.png
${DOC}kget/cr22-action-tool_queue.png
${DOC}kget/cr22-action-tool_restart.png
${DOC}kget/cr22-action-tool_resume.png
${DOC}kget/cr22-action-tool_shutdown.png
${DOC}kget/cr22-action-tool_timer.png
${DOC}kget/cr22-action-tool_uselastdir.png
${DOC}kget/${C}
${DOC}kget/${I}
${DOC}kget/kget1.png
${DOC}kget/kget2.png
${DOC}kget/kget3.png
${DOC}kget/kget4.png
${DOC}kget/kget5.png
${DOC}kghostview/common
${DOC}kghostview/${C}
${DOC}kghostview/${I}
${DOC}kgoldrunner/common
${DOC}kgoldrunner/editbar.png
${DOC}kgoldrunner/${C}
${DOC}kgoldrunner/${I}
${DOC}kgoldrunner/select.png
${DOC}kgoldrunner/tute008.png
${DOC}kgpg/common
${DOC}kgpg/editor.png
${DOC}kgpg/${C}
${DOC}kgpg/${I}
${DOC}kgpg/keygen.png
${DOC}kgpg/keymanage.png
${DOC}kgpg/keys.png
${DOC}kgpg/menu.png
${DOC}kgpg/options.png
${DOC}kgpgcertmanager/common
${DOC}kgpgcertmanager/${C}
${DOC}kgpgcertmanager/${I}
${DOC}khangman/common
${DOC}khangman/${C}
${DOC}khangman/${I}
${DOC}khangman/khangman1.png
${DOC}khangman/khangman2.png
${DOC}khelpcenter/common
${DOC}khelpcenter/contact.docbook
${DOC}khelpcenter/faq/about.docbook
${DOC}khelpcenter/faq/common
${DOC}khelpcenter/faq/configkde.docbook
${DOC}khelpcenter/faq/contrib.docbook
${DOC}khelpcenter/faq/desktop.docbook
${DOC}khelpcenter/faq/filemng.docbook
${DOC}khelpcenter/faq/getkde.docbook
${DOC}khelpcenter/faq/${C}
${DOC}khelpcenter/faq/${I}
${DOC}khelpcenter/faq/install.docbook
${DOC}khelpcenter/faq/intro.docbook
${DOC}khelpcenter/faq/kdeapps.docbook
${DOC}khelpcenter/faq/misc.docbook
${DOC}khelpcenter/faq/moreinfo.docbook
${DOC}khelpcenter/faq/nonkdeapps.docbook
${DOC}khelpcenter/faq/notrelated.docbook
${DOC}khelpcenter/faq/panel.docbook
${DOC}khelpcenter/faq/tips.docbook
${DOC}khelpcenter/faq/winmng.docbook
${DOC}khelpcenter/glossary/common
${DOC}khelpcenter/glossary/${C}
${DOC}khelpcenter/glossary/${I}
${DOC}khelpcenter/glossary/kdeprintingglossary.docbook
${DOC}khelpcenter/help.docbook
${DOC}khelpcenter/${C}
${DOC}khelpcenter/${I}
${DOC}khelpcenter/links.docbook
${DOC}khelpcenter/quickstart/common
${DOC}khelpcenter/quickstart/${C}
${DOC}khelpcenter/quickstart/${I}
${DOC}khelpcenter/support.docbook
${DOC}khelpcenter/userguide/about-desktop.docbook
${DOC}khelpcenter/userguide/common
${DOC}khelpcenter/userguide/first-impressions.docbook
${DOC}khelpcenter/userguide/getting-started.docbook
${DOC}khelpcenter/userguide/history.docbook
${DOC}khelpcenter/userguide/${C}
${DOC}khelpcenter/userguide/${I}
${DOC}khelpcenter/userguide/installation.docbook
${DOC}khelpcenter/userguide/intro.docbook
${DOC}khelpcenter/userguide/kdeadmin-apps.docbook
${DOC}khelpcenter/userguide/kdebase-apps.docbook
${DOC}khelpcenter/userguide/kdeedu-apps.docbook
${DOC}khelpcenter/userguide/kdegames-apps.docbook
${DOC}khelpcenter/userguide/kdegraphics-apps.docbook
${DOC}khelpcenter/userguide/kdemultimedia-apps.docbook
${DOC}khelpcenter/userguide/kdenetwork-apps.docbook
${DOC}khelpcenter/userguide/kdepim-apps.docbook
${DOC}khelpcenter/userguide/kdetoys-apps.docbook
${DOC}khelpcenter/userguide/kdeutils-apps.docbook
${DOC}khelpcenter/userguide/koffice-apps.docbook
${DOC}khelpcenter/userguide/more-help.docbook
${DOC}khelpcenter/userguide/notices-trademarks.docbook
${DOC}khelpcenter/userguide/shortcuts.docbook
${DOC}khelpcenter/userguide/staff.docbook
${DOC}khelpcenter/userguide/ug-faq.docbook
${DOC}khelpcenter/visualdict/common
${DOC}khelpcenter/visualdict/${C}
${DOC}khelpcenter/visualdict/${I}
${DOC}khelpcenter/welcome.docbook
${DOC}khelpcenter/whatiskde.docbook
${DOC}khexedit/common
${DOC}khexedit/${C}
${DOC}khexedit/${I}
${DOC}khexedit/khexedit1.png
${DOC}kicker-applets/common
${DOC}kicker-applets/${C}
${DOC}kicker-applets/${I}
${DOC}kicker-applets/kolourpicker.docbook
${DOC}kicker-applets/ktimemon.docbook
${DOC}kicker/common
${DOC}kicker/${C}
${DOC}kicker/${I}
${DOC}kiconedit/common
${DOC}kiconedit/${C}
${DOC}kiconedit/${I}
${DOC}kig/common
${DOC}kig/constructed_a_point.png
${DOC}kig/constructed_script_object.png
${DOC}kig/constructing_a_circle.png
${DOC}kig/constructing_a_circle_2.png
${DOC}kig/edit_types_dialog.png
${DOC}kig/${C}
${DOC}kig/${I}
${DOC}kig/macro_wizard.png
${DOC}kig/macros_at_work.png
${DOC}kig/script_wizard.png
${DOC}kig/script_wizard_entering_code.png
${DOC}kig/selecting_objects.png
${DOC}kig/simple_locus_construction.png
${DOC}kig/test_run_macro.png
${DOC}kig/text_label_attaching.png
${DOC}kig/text_label_wizard.png
${DOC}kig/text_label_wizard__select_property.png
${DOC}kinfocenter/blockdevices/common
${DOC}kinfocenter/blockdevices/${C}
${DOC}kinfocenter/blockdevices/${I}
${DOC}kinfocenter/common
${DOC}kinfocenter/devices/common
${DOC}kinfocenter/devices/${C}
${DOC}kinfocenter/devices/${I}
${DOC}kinfocenter/dma/common
${DOC}kinfocenter/dma/${C}
${DOC}kinfocenter/dma/${I}
${DOC}kinfocenter/${C}
${DOC}kinfocenter/${I}
${DOC}kinfocenter/interrupts/common
${DOC}kinfocenter/interrupts/${C}
${DOC}kinfocenter/interrupts/${I}
${DOC}kinfocenter/ioports/common
${DOC}kinfocenter/ioports/${C}
${DOC}kinfocenter/ioports/${I}
${DOC}kinfocenter/memory/common
${DOC}kinfocenter/memory/${C}
${DOC}kinfocenter/memory/${I}
${DOC}kinfocenter/nics/common
${DOC}kinfocenter/nics/${C}
${DOC}kinfocenter/nics/${I}
${DOC}kinfocenter/partitions/common
${DOC}kinfocenter/partitions/${C}
${DOC}kinfocenter/partitions/${I}
${DOC}kinfocenter/pci/common
${DOC}kinfocenter/pci/${C}
${DOC}kinfocenter/pci/${I}
${DOC}kinfocenter/pcmcia/common
${DOC}kinfocenter/pcmcia/${C}
${DOC}kinfocenter/pcmcia/${I}
${DOC}kinfocenter/processor/common
${DOC}kinfocenter/processor/${C}
${DOC}kinfocenter/processor/${I}
${DOC}kinfocenter/protocols/common
${DOC}kinfocenter/protocols/${C}
${DOC}kinfocenter/protocols/${I}
${DOC}kinfocenter/samba/common
${DOC}kinfocenter/samba/${C}
${DOC}kinfocenter/samba/${I}
${DOC}kinfocenter/scsi/common
${DOC}kinfocenter/scsi/${C}
${DOC}kinfocenter/scsi/${I}
${DOC}kinfocenter/sound/common
${DOC}kinfocenter/sound/${C}
${DOC}kinfocenter/sound/${I}
${DOC}kinfocenter/usb/common
${DOC}kinfocenter/usb/${C}
${DOC}kinfocenter/usb/${I}
${DOC}kinfocenter/xserver/common
${DOC}kinfocenter/xserver/${C}
${DOC}kinfocenter/xserver/${I}
${DOC}kioslave/audiocd.docbook
${DOC}kioslave/bzip.docbook
${DOC}kioslave/bzip2.docbook
${DOC}kioslave/cgi.docbook
${DOC}kioslave/common
${DOC}kioslave/data.docbook
${DOC}kioslave/file.docbook
${DOC}kioslave/finger.docbook
${DOC}kioslave/fish.docbook
${DOC}kioslave/floppy.docbook
${DOC}kioslave/ftp.docbook
${DOC}kioslave/gopher.docbook
${DOC}kioslave/gzip.docbook
${DOC}kioslave/help.docbook
${DOC}kioslave/http.docbook
${DOC}kioslave/https.docbook
${DOC}kioslave/imap.docbook
${DOC}kioslave/imaps.docbook
${DOC}kioslave/${C}
${DOC}kioslave/${I}
${DOC}kioslave/info.docbook
${DOC}kioslave/lan.docbook
${DOC}kioslave/ldap.docbook
${DOC}kioslave/mac.docbook
${DOC}kioslave/mailto.docbook
${DOC}kioslave/man.docbook
${DOC}kioslave/mrml.docbook
${DOC}kioslave/news.docbook
${DOC}kioslave/nfs.docbook
${DOC}kioslave/nntp.docbook
${DOC}kioslave/pop3.docbook
${DOC}kioslave/pop3s.docbook
${DOC}kioslave/print.docbook
${DOC}kioslave/rdate.docbook
${DOC}kioslave/rlan.docbook
${DOC}kioslave/rlogin.docbook
${DOC}kioslave/sftp.docbook
${DOC}kioslave/smb.docbook
${DOC}kioslave/smtp.docbook
${DOC}kioslave/tar.docbook
${DOC}kioslave/telnet.docbook
${DOC}kioslave/thumbnail.docbook
${DOC}kioslave/webdav.docbook
${DOC}kioslave/webdavs.docbook
${DOC}kit/common
${DOC}kit/${C}
${DOC}kit/${I}
${DOC}kiten/common
${DOC}kiten/${C}
${DOC}kiten/${I}
${DOC}kjots/common
${DOC}kjots/${C}
${DOC}kjots/${I}
${DOC}kjumpingcube/common
${DOC}kjumpingcube/${C}
${DOC}kjumpingcube/${I}
${DOC}klettres/common
${DOC}klettres/${C}
${DOC}klettres/${I}
${DOC}klettres/klettres1.png
${DOC}klettres/klettres2.png
${DOC}klettres/klettres3.png
${DOC}klettres/klettres4.png
${DOC}klettres/klettres5.png
${DOC}klickety/common
${DOC}klickety/${C}
${DOC}klickety/${I}
${DOC}klines/common
${DOC}klines/${C}
${DOC}klines/${I}
${DOC}klipper/common
${DOC}klipper/${C}
${DOC}klipper/${I}
${DOC}kmag/common
${DOC}kmag/images/screenshot.png
${DOC}kmag/${C}
${DOC}kmag/${I}
${DOC}kmag/screenshot.png
${DOC}kmail/common
${DOC}kmail/configure.docbook
${DOC}kmail/credits-and-licenses.docbook
${DOC}kmail/faq.docbook
${DOC}kmail/getting-started.docbook
${DOC}kmail/importing.docbook
${DOC}kmail/${C}
${DOC}kmail/${I}
${DOC}kmail/intro.docbook
${DOC}kmail/menus.docbook
${DOC}kmail/using-kmail.docbook
${DOC}kmathtool/common
${DOC}kmathtool/${C}
${DOC}kmathtool/${I}
${DOC}kmenuedit/common
${DOC}kmenuedit/${C}
${DOC}kmenuedit/${I}
${DOC}kmessedwords/common
${DOC}kmessedwords/${C}
${DOC}kmessedwords/${I}
${DOC}kmessedwords/kmw1.png
${DOC}kmessedwords/kmw2.png
${DOC}kmessedwords/kmw3.png
${DOC}kmessedwords/kmw4.png
${DOC}kmid/common
${DOC}kmid/${C}
${DOC}kmid/${I}
${DOC}kmidi/common
${DOC}kmidi/${C}
${DOC}kmidi/${I}
${DOC}kmines/common
${DOC}kmines/${C}
${DOC}kmines/${I}
${DOC}kmines/kmines1.png
${DOC}kmines/kmines2.png
${DOC}kmix/common
${DOC}kmix/${C}
${DOC}kmix/${I}
${DOC}kmoon/common
${DOC}kmoon/${C}
${DOC}kmoon/${I}
${DOC}kmousetool/common
${DOC}kmousetool/${C}
${DOC}kmousetool/${I}
${DOC}kmouth/common
${DOC}kmouth/${C}
${DOC}kmouth/${I}
${DOC}kmouth/kmouthctts.png
${DOC}kmouth/kmouthedit.png
${DOC}kmouth/kmouthmain.png
${DOC}kmouth/kmouthwizard.png
${DOC}kmplot/commands.docbook
${DOC}kmplot/common
${DOC}kmplot/configuration.docbook
${DOC}kmplot/credits.docbook
${DOC}kmplot/developer.docbook
${DOC}kmplot/${C}
${DOC}kmplot/${I}
${DOC}kmplot/install.docbook
${DOC}kmplot/introduction.docbook
${DOC}kmplot/main.png
${DOC}kmplot/menu.docbook
${DOC}kmplot/namesdlg.png
${DOC}kmplot/reference.docbook
${DOC}kmplot/using.docbook
${DOC}knewsticker/common
${DOC}knewsticker/contextmenu.png
${DOC}knewsticker/${C}
${DOC}knewsticker/${I}
${DOC}knewsticker/kcmnewsticker-filters.png
${DOC}knewsticker/kcmnewsticker-general.png
${DOC}knewsticker/kcmnewsticker-newssitedialog.png
${DOC}knewsticker/kcmnewsticker-newssources.png
${DOC}knewsticker/kcmnewsticker-scrollerprefs.png
${DOC}knode/commands.docbook
${DOC}knode/common
${DOC}knode/credits.docbook
${DOC}knode/faq.docbook
${DOC}knode/gloss.docbook
${DOC}knode/${C}
${DOC}knode/${I}
${DOC}knode/install.docbook
${DOC}knode/introduction.docbook
${DOC}knode/journey.docbook
${DOC}knode/knode-cleanup.png
${DOC}knode/knode-colors-fonts.png
${DOC}knode/knode-composer-attachments.png
${DOC}knode/knode-composer-settings.png
${DOC}knode/knode-edit-filter.png
${DOC}knode/knode-edit-header1.png
${DOC}knode/knode-edit-header2.png
${DOC}knode/knode-filters.png
${DOC}knode/knode-followup.png
${DOC}knode/knode-header-settings.png
${DOC}knode/knode-identity.png
${DOC}knode/knode-mail-account.png
${DOC}knode/knode-new-article.png
${DOC}knode/knode-news-account.png
${DOC}knode/knode-post-settings.png
${DOC}knode/knode-read-news-settings.png
${DOC}knode/knode-reply.png
${DOC}knode/knode-rule-editor.png
${DOC}knode/knode-search.png
${DOC}knode/knode-start.png
${DOC}knode/knode-subscribe.png
${DOC}knode/knode-views.png
${DOC}knode/more.docbook
${DOC}knode/using-firststart.docbook
${DOC}knode/using-morefeatures.docbook
${DOC}knode/using-subscribing.docbook
${DOC}knotes/common
${DOC}knotes/${C}
${DOC}knotes/${I}
${DOC}kodo/common
${DOC}kodo/${C}
${DOC}kodo/${I}
${DOC}kolf/common
${DOC}kolf/${C}
${DOC}kolf/${I}
${DOC}kompare/common
${DOC}kompare/${C}
${DOC}kompare/${I}
${DOC}konq-plugins/babel/common
${DOC}konq-plugins/babel/${C}
${DOC}konq-plugins/babel/${I}
${DOC}konq-plugins/common
${DOC}konq-plugins/crashes/common
${DOC}konq-plugins/crashes/${C}
${DOC}konq-plugins/crashes/${I}
${DOC}konq-plugins/dirfilter/common
${DOC}konq-plugins/dirfilter/${C}
${DOC}konq-plugins/dirfilter/${I}
${DOC}konq-plugins/domtreeviewer/common
${DOC}konq-plugins/domtreeviewer/${C}
${DOC}konq-plugins/domtreeviewer/${I}
${DOC}konq-plugins/fsview/common
${DOC}konq-plugins/fsview/${C}
${DOC}konq-plugins/fsview/${I}
${DOC}konq-plugins/imgallery/common
${DOC}konq-plugins/imgallery/${C}
${DOC}konq-plugins/imgallery/${I}
${DOC}konq-plugins/${C}
${DOC}konq-plugins/${I}
${DOC}konq-plugins/khtmlsettings/common
${DOC}konq-plugins/khtmlsettings/${C}
${DOC}konq-plugins/khtmlsettings/${I}
${DOC}konq-plugins/kuick/common
${DOC}konq-plugins/kuick/${C}
${DOC}konq-plugins/kuick/${I}
${DOC}konq-plugins/mediaplayer/common
${DOC}konq-plugins/mediaplayer/${C}
${DOC}konq-plugins/mediaplayer/${I}
${DOC}konq-plugins/smbmounter/common
${DOC}konq-plugins/smbmounter/${C}
${DOC}konq-plugins/smbmounter/${I}
${DOC}konq-plugins/uachanger/common
${DOC}konq-plugins/uachanger/${C}
${DOC}konq-plugins/uachanger/${I}
${DOC}konq-plugins/validators/common
${DOC}konq-plugins/validators/${C}
${DOC}konq-plugins/validators/${I}
${DOC}konq-plugins/webarchiver/common
${DOC}konq-plugins/webarchiver/${C}
${DOC}konq-plugins/webarchiver/${I}
${DOC}konqueror/basics.docbook
${DOC}konqueror/bookmarks.docbook
${DOC}konqueror/browser.docbook
${DOC}konqueror/cmndline.png
${DOC}konqueror/commands.docbook
${DOC}konqueror/common
${DOC}konqueror/config.docbook
${DOC}konqueror/credits.docbook
${DOC}konqueror/dirtree.png
${DOC}konqueror/dragdrop.png
${DOC}konqueror/faq.docbook
${DOC}konqueror/filemanager.docbook
${DOC}konqueror/filetype1.png
${DOC}konqueror/filetype3.png
${DOC}konqueror/filetype4.png
${DOC}konqueror/${C}
${DOC}konqueror/${I}
${DOC}konqueror/introduction.docbook
${DOC}konqueror/konqorg.png
${DOC}konqueror/parts.png
${DOC}konqueror/path-complete.docbook
${DOC}konqueror/plugins.docbook
${DOC}konqueror/save-settings.docbook
${DOC}konqueror/shortcut1.png
${DOC}konqueror/shortcut2.png
${DOC}konqueror/sidebar.docbook
${DOC}konquest/common
${DOC}konquest/${C}
${DOC}konquest/${I}
${DOC}konsole/common
${DOC}konsole/${C}
${DOC}konsole/${I}
${DOC}konsole/konsole.png
${DOC}konsolekalendar/common
${DOC}konsolekalendar/${C}
${DOC}konsolekalendar/${I}
${DOC}kontact/common
${DOC}kontact/${C}
${DOC}kontact/${I}
${DOC}kooka/common
${DOC}kooka/${C}
${DOC}kooka/${I}
${DOC}kooka/kooka_gocr.png
${DOC}kooka/kooka_gocr_result.png
${DOC}kooka/kooka_mainctrl.png
${DOC}kooka/shortcut0.png
${DOC}kooka/shortcut1.png
${DOC}kooka/toolbar.png
${DOC}kooka/toolbar1.png
${DOC}kooka/toolbar2.png
${DOC}kopete/common
${DOC}kopete/${C}
${DOC}kopete/${I}
${DOC}korganizer/common
${DOC}korganizer/ep_config.png
${DOC}korganizer/ep_download.png
${DOC}korganizer/ep_enable.png
${DOC}korganizer/ep_menu.png
${DOC}korganizer/ep_progress.png
${DOC}korganizer/exchange-plugin.docbook
${DOC}korganizer/group-scheduling.docbook
${DOC}korganizer/gs_attendee1.png
${DOC}korganizer/gs_attendee2.png
${DOC}korganizer/gs_counter.png
${DOC}korganizer/gs_filter.png
${DOC}korganizer/gs_inbox1.png
${DOC}korganizer/gs_inbox2.png
${DOC}korganizer/gs_korganizer1.png
${DOC}korganizer/gs_korganizer2.png
${DOC}korganizer/gs_korganizer3.png
${DOC}korganizer/gs_outbox1.png
${DOC}korganizer/gs_outbox2.png
${DOC}korganizer/gs_publish.png
${DOC}korganizer/gs_reply.png
${DOC}korganizer/gs_setup1.png
${DOC}korganizer/gs_setup2.png
${DOC}korganizer/gs_show1.png
${DOC}korganizer/gs_show2.png
${DOC}korganizer/gs_whatsnext.png
${DOC}korganizer/${C}
${DOC}korganizer/${I}
${DOC}korganizer/o2v_importing1.png
${DOC}korganizer/o2v_importing2.png
${DOC}korganizer/o2v_importing3.png
${DOC}korganizer/outlook-to-vcalendar.docbook
${DOC}korn/common
${DOC}korn/${C}
${DOC}korn/${I}
${DOC}kpackage/bsdloc.png
${DOC}kpackage/common
${DOC}kpackage/debaptloc.png
${DOC}kpackage/debloc.png
${DOC}kpackage/handle.png
${DOC}kpackage/${C}
${DOC}kpackage/${I}
${DOC}kpackage/install.png
${DOC}kpackage/left.png
${DOC}kpackage/right-change.png
${DOC}kpackage/right-files.png
${DOC}kpackage/right-prop.png
${DOC}kpackage/rpmloc.png
${DOC}kpackage/slackloc.png
${DOC}kpackage/uninstall.png
${DOC}kpager/common
${DOC}kpager/${C}
${DOC}kpager/${I}
${DOC}kpager/screenshot.png
${DOC}kpager/settings.png
${DOC}kpaint/common
${DOC}kpaint/${C}
${DOC}kpaint/${I}
${DOC}kpat/common
${DOC}kpat/${C}
${DOC}kpat/${I}
${DOC}kpat/man.docbook
${DOC}kpdf/common
${DOC}kpdf/${C}
${DOC}kpdf/${I}
${DOC}kpercentage/answer.png
${DOC}kpercentage/commands.docbook
${DOC}kpercentage/common
${DOC}kpercentage/credits.docbook
${DOC}kpercentage/devel.docbook
${DOC}kpercentage/faq.docbook
${DOC}kpercentage/help.png
${DOC}kpercentage/${C}
${DOC}kpercentage/${I}
${DOC}kpercentage/install.docbook
${DOC}kpercentage/introduction.docbook
${DOC}kpercentage/main.png
${DOC}kpercentage/using.docbook
${DOC}kpercentage/welcome.png
${DOC}kpf/common
${DOC}kpf/${C}
${DOC}kpf/${I}
${DOC}kpilot/address-app.png
${DOC}kpilot/common
${DOC}kpilot/conduit-knotes.png
${DOC}kpilot/conduit-popmail-kmail.png
${DOC}kpilot/conduit-popmail-recv-method.png
${DOC}kpilot/conduit-popmail-send-as.png
${DOC}kpilot/conduit-popmail-send-method.png
${DOC}kpilot/conduit-popmail-sendmail.png
${DOC}kpilot/conduit-popmail-smtp.png
${DOC}kpilot/conduit-popmail-top.png
${DOC}kpilot/conduit-vcal.png
${DOC}kpilot/file-app.png
${DOC}kpilot/${C}
${DOC}kpilot/${I}
${DOC}kpilot/main-app.png
${DOC}kpilot/memo-app.png
${DOC}kpilot/setup-address.png
${DOC}kpilot/setup-conduit.png
${DOC}kpilot/setup-dbspecial.png
${DOC}kpilot/setup-general.png
${DOC}kpilot/setup-sync.png
${DOC}kpoker/common
${DOC}kpoker/${C}
${DOC}kpoker/${I}
${DOC}kpoker/kpoker1.png
${DOC}kpoker/kpoker2.png
${DOC}kpovmodeler/cameraview.png
${DOC}kpovmodeler/common
${DOC}kpovmodeler/controlpoints.png
${DOC}kpovmodeler/defaultviewlayout.png
${DOC}kpovmodeler/dockwidget.png
${DOC}kpovmodeler/dockwidgettab.png
${DOC}kpovmodeler/${C}
${DOC}kpovmodeler/${I}
${DOC}kpovmodeler/insertaspopup.png
${DOC}kpovmodeler/objectpropertiesview.png
${DOC}kpovmodeler/objecttree.png
${DOC}kpovmodeler/rendermodeoutput.png
${DOC}kpovmodeler/rendermodequality.png
${DOC}kpovmodeler/rendermodesize.png
${DOC}kpovmodeler/rendermodesselection.png
${DOC}kpovmodeler/rendermodestoolbar.png
${DOC}kpovmodeler/renderwindow.png
${DOC}kpovmodeler/texturepreview.png
${DOC}kpovmodeler/topview.png
${DOC}kpovmodeler/tutorial01-camera-dialog.png
${DOC}kpovmodeler/tutorial01-camera-graphic.png
${DOC}kpovmodeler/tutorial01-ground-color-list.png
${DOC}kpovmodeler/tutorial01-ground-pigment.png
${DOC}kpovmodeler/tutorial01-ground-render.png
${DOC}kpovmodeler/tutorial01-ground-solid-color-1.png
${DOC}kpovmodeler/tutorial01-ground-solid-color-2.png
${DOC}kpovmodeler/tutorial01-ground-wrong-colors-render.png
${DOC}kpovmodeler/tutorial01-light-dialog.png
${DOC}kpovmodeler/tutorial01-light-graphic.png
${DOC}kpovmodeler/tutorial01-plane-dialog.png
${DOC}kpovmodeler/tutorial01-plane-graphic.png
${DOC}kpovmodeler/tutorial01-plane-tree-expanded.png
${DOC}kpovmodeler/tutorial01-plane-tree-translate.png
${DOC}kpovmodeler/tutorial01-sphere-dialog.png
${DOC}kpovmodeler/tutorial01-sphere-finish-dialog.png
${DOC}kpovmodeler/tutorial01-sphere-render-finish.png
${DOC}kpovmodeler/tutorial01-sphere-render-nocolor.png
${DOC}kpovmodeler/tutorial01-sphere-render-solidcolor.png
${DOC}kpovmodeler/tutorial01-sphere-solid-color.png
${DOC}kppp/accounting.docbook
${DOC}kppp/callback.docbook
${DOC}kppp/chap.docbook
${DOC}kppp/common
${DOC}kppp/dialog-setup.docbook
${DOC}kppp/getting-online.docbook
${DOC}kppp/global-settings.docbook
${DOC}kppp/hayes.docbook
${DOC}kppp/${C}
${DOC}kppp/${I}
${DOC}kppp/kppp-account-accounting-tab.png
${DOC}kppp/kppp-account-dial-tab.png
${DOC}kppp/kppp-account-dns-tab.png
${DOC}kppp/kppp-account-execute-tab.png
${DOC}kppp/kppp-account-gateway-tab.png
${DOC}kppp/kppp-account-ip-tab.png
${DOC}kppp/kppp-account-login-script-tab.png
${DOC}kppp/kppp-config.png
${DOC}kppp/kppp-device-tab.png
${DOC}kppp/kppp-dialler-tab.png
${DOC}kppp/kppp-faq.docbook
${DOC}kppp/kppp-graph-tab.png
${DOC}kppp/kppp-misc-tab.png
${DOC}kppp/kppp-modem-tab.png
${DOC}kppp/kppp-wizard.png
${DOC}kppp/security.docbook
${DOC}kppp/tricks.docbook
${DOC}kppp/wizard.docbook
${DOC}krdc/authentication.png
${DOC}krdc/common
${DOC}krdc/${C}
${DOC}krdc/${I}
${DOC}krdc/preferences_profilestab.png
${DOC}krdc/preferences_rdpdefaultstab.png
${DOC}krdc/preferences_vncdefaultstab.png
${DOC}krdc/snapshot.png
${DOC}krdc/snapshot_connectionspeed.png
${DOC}krdc/snapshot_nobrowse.png
${DOC}krdc/snapshot_vncentry.png
${DOC}krec/common
${DOC}krec/${C}
${DOC}krec/${I}
${DOC}krec/krec-hicolor.png
${DOC}kreversi/common
${DOC}kreversi/${C}
${DOC}kreversi/${I}
${DOC}kreversi/kreversi1.png
${DOC}krfb/common
${DOC}krfb/configuration_access.png
${DOC}krfb/configuration_network.png
${DOC}krfb/configuration_session.png
${DOC}krfb/connection.png
${DOC}krfb/email_invitation.png
${DOC}krfb/${C}
${DOC}krfb/${I}
${DOC}krfb/invitation_management.png
${DOC}krfb/personal_invitation.png
${DOC}krfb/screenshot.png
${DOC}kruler/common
${DOC}kruler/${C}
${DOC}kruler/${I}
${DOC}ksame/common
${DOC}ksame/${C}
${DOC}ksame/${I}
${DOC}kscd/common
${DOC}kscd/${C}
${DOC}kscd/${I}
${DOC}kscd/kscd.png
${DOC}kscd/kscd12.png
${DOC}kscd/kscd13.png
${DOC}kscd/kscd14.png
${DOC}kscd/kscd16.png
${DOC}kscd/kscd19.png
${DOC}kscd/kscd2.png
${DOC}kscd/kscd3.png
${DOC}kshisen/common
${DOC}kshisen/${C}
${DOC}kshisen/${I}
${DOC}ksim/common
${DOC}ksim/${C}
${DOC}ksim/${I}
${DOC}ksirc/common
${DOC}ksirc/${C}
${DOC}ksirc/${I}
${DOC}ksirtet/common
${DOC}ksirtet/${C}
${DOC}ksirtet/${I}
${DOC}ksnake/common
${DOC}ksnake/${C}
${DOC}ksnake/${I}
${DOC}ksnapshot/common
${DOC}ksnapshot/${C}
${DOC}ksnapshot/${I}
${DOC}ksnapshot/preview.png
${DOC}ksnapshot/window.png
${DOC}ksokoban/common
${DOC}ksokoban/${C}
${DOC}ksokoban/${I}
${DOC}kspaceduel/common
${DOC}kspaceduel/${C}
${DOC}kspaceduel/${I}
${DOC}kspaceduel/kspaceduel1.png
${DOC}kspaceduel/kspaceduel2.png
${DOC}kspaceduel/kspaceduel3.png
${DOC}kspell/common
${DOC}kspell/${C}
${DOC}kspell/${I}
${DOC}ksplashml/common
${DOC}ksplashml/${C}
${DOC}ksplashml/${I}
${DOC}kstars/aavso.png
${DOC}kstars/ai-contents.docbook
${DOC}kstars/altvstime.docbook
${DOC}kstars/altvstime.png
${DOC}kstars/astroinfo.docbook
${DOC}kstars/blackbody.docbook
${DOC}kstars/blackbody.png
${DOC}kstars/calc-apcoords.docbook
${DOC}kstars/calc-apcoords.png
${DOC}kstars/calc-dayduration.docbook
${DOC}kstars/calc-daylength.png
${DOC}kstars/calc-eqgal.docbook
${DOC}kstars/calc-eqgal.png
${DOC}kstars/calc-geodetic.docbook
${DOC}kstars/calc-geodetic.png
${DOC}kstars/calc-horizontal.docbook
${DOC}kstars/calc-horizontal.png
${DOC}kstars/calc-julian.png
${DOC}kstars/calc-julianday.docbook
${DOC}kstars/calc-precess.docbook
${DOC}kstars/calc-precess.png
${DOC}kstars/calc-sidereal.docbook
${DOC}kstars/calc-sidereal.png
${DOC}kstars/calculator.docbook
${DOC}kstars/cequator.docbook
${DOC}kstars/color_indices.png
${DOC}kstars/colorandtemp.docbook
${DOC}kstars/commands.docbook
${DOC}kstars/common
${DOC}kstars/config.docbook
${DOC}kstars/cpoles.docbook
${DOC}kstars/credits.docbook
${DOC}kstars/csphere.docbook
${DOC}kstars/darkmatter.docbook
${DOC}kstars/dcop.docbook
${DOC}kstars/detaildialog.png
${DOC}kstars/details.docbook
${DOC}kstars/devicemanager.png
${DOC}kstars/dumpmode.docbook
${DOC}kstars/ecliptic.docbook
${DOC}kstars/ellipticalgalaxies.docbook
${DOC}kstars/equinox.docbook
${DOC}kstars/faq.docbook
${DOC}kstars/find.png
${DOC}kstars/flux.docbook
${DOC}kstars/fovdialog.png
${DOC}kstars/geocoords.docbook
${DOC}kstars/geolocator.png
${DOC}kstars/greatcircle.docbook
${DOC}kstars/horizon.docbook
${DOC}kstars/hourangle.docbook
${DOC}kstars/${C}
${DOC}kstars/${I}
${DOC}kstars/indi.docbook
${DOC}kstars/indiclient.png
${DOC}kstars/indicontrolpanel.png
${DOC}kstars/install.docbook
${DOC}kstars/jmoons.docbook
${DOC}kstars/jmoons.png
${DOC}kstars/julianday.docbook
${DOC}kstars/leapyear.docbook
${DOC}kstars/lightcurve.png
${DOC}kstars/lightcurves.docbook
${DOC}kstars/luminosity.docbook
${DOC}kstars/magnitude.docbook
${DOC}kstars/meridian.docbook
${DOC}kstars/newfov.png
${DOC}kstars/parallax.docbook
${DOC}kstars/popup.png
${DOC}kstars/precession.docbook
${DOC}kstars/quicktour.docbook
${DOC}kstars/retrograde.docbook
${DOC}kstars/screen1.png
${DOC}kstars/scriptbuilder.docbook
${DOC}kstars/scriptbuilder.png
${DOC}kstars/sidereal.docbook
${DOC}kstars/skycoords.docbook
${DOC}kstars/skymapdevice.png
${DOC}kstars/solarsys.docbook
${DOC}kstars/solarsystem.png
${DOC}kstars/spiralgalaxies.docbook
${DOC}kstars/star_colors.png
${DOC}kstars/stars.docbook
${DOC}kstars/timezones.docbook
${DOC}kstars/tools.docbook
${DOC}kstars/utime.docbook
${DOC}kstars/viewops.png
${DOC}kstars/wut.docbook
${DOC}kstars/wut.png
${DOC}kstars/zenith.docbook
${DOC}ksysguard/common
${DOC}ksysguard/${C}
${DOC}ksysguard/${I}
${DOC}ksysv/common
${DOC}ksysv/${C}
${DOC}ksysv/${I}
${DOC}ktalkd/common
${DOC}ktalkd/${C}
${DOC}ktalkd/${I}
${DOC}kteatime/common
${DOC}kteatime/config.png
${DOC}kteatime/${C}
${DOC}kteatime/${I}
${DOC}ktimer/common
${DOC}ktimer/${C}
${DOC}ktimer/${I}
${DOC}ktouch/common
${DOC}ktouch/${C}
${DOC}ktouch/${I}
${DOC}ktouch/screenshot1.png
${DOC}ktouch/screenshot2.png
${DOC}ktouch/screenshot3.png
${DOC}ktron/common
${DOC}ktron/${C}
${DOC}ktron/${I}
${DOC}ktuberling/common
${DOC}ktuberling/${C}
${DOC}ktuberling/${I}
${DOC}ktuberling/menu.edit.png
${DOC}ktuberling/menu.file.png
${DOC}ktuberling/menu.game.png
${DOC}ktuberling/menu.help.png
${DOC}ktuberling/menu.option.png
${DOC}ktuberling/menu.playground.png
${DOC}ktuberling/menu.raw.png
${DOC}ktuberling/menu.speech.png
${DOC}ktuberling/technical-reference.docbook
${DOC}kuickshow/common
${DOC}kuickshow/${C}
${DOC}kuickshow/${I}
${DOC}kuickshow/screenshot.png
${DOC}kuser/common
${DOC}kuser/${C}
${DOC}kuser/${I}
${DOC}kverbos/common
${DOC}kverbos/${C}
${DOC}kverbos/${I}
${DOC}kverbos/input.png
${DOC}kverbos/mainscreen-leer.png
${DOC}kverbos/mainscreen1.png
${DOC}kverbos/newverb.png
${DOC}kverbos/options.png
${DOC}kverbos/result.png
${DOC}kverbos/type.png
${DOC}kverbos/username.png
${DOC}kverbos/verblist.png
${DOC}kview/common
${DOC}kview/${C}
${DOC}kview/${I}
${DOC}kview/snapshot1.png
${DOC}kview/snapshot2.png
${DOC}kview/snapshot3.png
${DOC}kview/snapshot4.png
${DOC}kview/snapshot5.png
${DOC}kview/snapshot6.png
${DOC}kview/snapshot7.png
${DOC}kview/snapshot8.png
${DOC}kview/snapshot9.png
${DOC}kvoctrain/art-query-dlg.png
${DOC}kvoctrain/common
${DOC}kvoctrain/comp-query-dlg.png
${DOC}kvoctrain/docprop1-dlg.png
${DOC}kvoctrain/docprop2-dlg.png
${DOC}kvoctrain/docprop6-dlg.png
${DOC}kvoctrain/entry1-dlg.png
${DOC}kvoctrain/entry2-dlg.png
${DOC}kvoctrain/entry3-dlg.png
${DOC}kvoctrain/entry4-dlg.png
${DOC}kvoctrain/entry5-dlg.png
${DOC}kvoctrain/entry6-dlg.png
${DOC}kvoctrain/${C}
${DOC}kvoctrain/${I}
${DOC}kvoctrain/lang1-dlg.png
${DOC}kvoctrain/mainview.png
${DOC}kvoctrain/mu-query-dlg.png
${DOC}kvoctrain/options1-dlg.png
${DOC}kvoctrain/options2-dlg.png
${DOC}kvoctrain/options3-dlg.png
${DOC}kvoctrain/options4-dlg.png
${DOC}kvoctrain/pron-dlg.png
${DOC}kvoctrain/q-opt1-dlg.png
${DOC}kvoctrain/q-opt2-dlg.png
${DOC}kvoctrain/q-opt3-dlg.png
${DOC}kvoctrain/q-opt4-dlg.png
${DOC}kvoctrain/query-dlg.png
${DOC}kvoctrain/stat1-dlg.png
${DOC}kvoctrain/stat2-dlg.png
${DOC}kvoctrain/syn-query-dlg.png
${DOC}kvoctrain/verb-query-dlg.png
${DOC}kwallet/common
${DOC}kwallet/${C}
${DOC}kwallet/${I}
${DOC}kweather/common
${DOC}kweather/${C}
${DOC}kweather/${I}
${DOC}kwifimanager/common
${DOC}kwifimanager/${C}
${DOC}kwifimanager/${I}
${DOC}kwin4/common
${DOC}kwin4/${C}
${DOC}kwin4/${I}
${DOC}kworldclock/common
${DOC}kworldclock/${C}
${DOC}kworldclock/${I}
${DOC}kwrite/common
${DOC}kwrite/${C}
${DOC}kwrite/${I}
${DOC}kwuftpd/common
${DOC}kwuftpd/directories.png
${DOC}kwuftpd/${C}
${DOC}kwuftpd/${I}
${DOC}kwuftpd/logging.png
${DOC}kwuftpd/messages.png
${DOC}kwuftpd/ratios.png
${DOC}kwuftpd/security.png
${DOC}kwuftpd/uploads.png
${DOC}kwuftpd/user_classes.png
${DOC}kwuftpd/virtual.png
${DOC}kxconfig/common
${DOC}kxconfig/${C}
${DOC}kxconfig/${I}
${DOC}kxkb/common
${DOC}kxkb/${C}
${DOC}kxkb/${I}
${DOC}kxsldbg/breakpoints_window.png
${DOC}kxsldbg/callstack.docbook
${DOC}kxsldbg/callstack_window.png
${DOC}kxsldbg/common
${DOC}kxsldbg/configure_window.png
${DOC}kxsldbg/credits.docbook
${DOC}kxsldbg/entities.docbook
${DOC}kxsldbg/entities_window.png
${DOC}kxsldbg/globals_window.png
${DOC}kxsldbg/glossary.docbook
${DOC}kxsldbg/${C}
${DOC}kxsldbg/${I}
${DOC}kxsldbg/kxsldbg_configure.docbook
${DOC}kxsldbg/kxsldbg_inspector.docbook
${DOC}kxsldbg/kxsldbg_mainwindow.docbook
${DOC}kxsldbg/kxsldbg_tools.docbook
${DOC}kxsldbg/main_window.png
${DOC}kxsldbg/publicid_window.png
${DOC}kxsldbg/sources.docbook
${DOC}kxsldbg/sources_window.png
${DOC}kxsldbg/systemid_window.png
${DOC}kxsldbg/templates.docbook
${DOC}kxsldbg/templates_window.png
${DOC}kxsldbg/variables.docbook
${DOC}kxsldbg/walk_window.png
${DOC}lisa/common
${DOC}lisa/${C}
${DOC}lisa/${I}
${DOC}lskat/common
${DOC}lskat/${C}
${DOC}lskat/${I}
${DOC}megami/common
${DOC}megami/${C}
${DOC}megami/${I}
${DOC}noatun/common
${DOC}noatun/${C}
${DOC}noatun/${I}
${DOC}quanta/adv-quanta.docbook
${DOC}quanta/attribute_tree.png
${DOC}quanta/common
${DOC}quanta/conf-action.png
${DOC}quanta/conf-action1.png
${DOC}quanta/conf-action2.png
${DOC}quanta/config-quanta.docbook
${DOC}quanta/credits-license.docbook
${DOC}quanta/debugging-quanta.docbook
${DOC}quanta/doc-view1.png
${DOC}quanta/dtep_doc_img15.png
${DOC}quanta/dtep_doc_img18.png
${DOC}quanta/dtep_doc_img21.png
${DOC}quanta/dtep_doc_img22.png
${DOC}quanta/dtep_doc_img23.png
${DOC}quanta/dtep_doc_img24.png
${DOC}quanta/dtep_doc_img25.png
${DOC}quanta/dtep_doc_img7.png
${DOC}quanta/dtep_doc_img8.png
${DOC}quanta/extending-quanta.docbook
${DOC}quanta/fundamentals.docbook
${DOC}quanta/glossary.docbook
${DOC}quanta/${C}
${DOC}quanta/${I}
${DOC}quanta/installation.docbook
${DOC}quanta/introduction.docbook
${DOC}quanta/plugin-edit.png
${DOC}quanta/project-1.png
${DOC}quanta/project-tree-view-dir-rmb-menu.png
${DOC}quanta/project-tree-view-file-rmb-menu.png
${DOC}quanta/project-upload-dialog.png
${DOC}quanta/q-and-a.docbook
${DOC}quanta/quanta-menus.docbook
${DOC}quanta/quanta-projects.docbook
${DOC}quanta/quantamdi-editor.png
${DOC}quanta/quantamdi-treeview.png
${DOC}quanta/quantamdi.png
${DOC}quanta/taginputex.png
${DOC}quanta/template-rmb.png
${DOC}quanta/toolbars.png
${DOC}quanta/using-quanta.docbook
${DOC}quanta/vplsourceview.png
${DOC}quanta/working-with-quanta.docbook
${DOC}umbrello/authors.docbook
${DOC}umbrello/code_import_and_generation.docbook
${DOC}umbrello/common
${DOC}umbrello/credits.docbook
${DOC}umbrello/faq.docbook
${DOC}umbrello/${C}
${DOC}umbrello/${I}
${DOC}umbrello/installation.docbook
${DOC}umbrello/introduction.docbook
${DOC}umbrello/other_features.docbook
${DOC}umbrello/pics/activity-diagram.png
${DOC}umbrello/pics/add-remove-languages.png
${DOC}umbrello/pics/aggregation.png
${DOC}umbrello/pics/association.png
${DOC}umbrello/pics/class-diagram.png
${DOC}umbrello/pics/class.png
${DOC}umbrello/pics/code-import.png
${DOC}umbrello/pics/collaboration-diagram.png
${DOC}umbrello/pics/composition.png
${DOC}umbrello/pics/folders.png
${DOC}umbrello/pics/generalization.png
${DOC}umbrello/pics/generation-options.png
${DOC}umbrello/pics/sequence-diagram.png
${DOC}umbrello/pics/state-diagram.png
${DOC}umbrello/pics/umbrello-main-screen.png
${DOC}umbrello/pics/umbrello-ui.png
${DOC}umbrello/pics/use-case-diagram.png
${DOC}umbrello/uml_basics.docbook
${DOC}umbrello/working_with_umbrello.docbook
${LOC}alarmdaemonctrl.mo
${LOC}alsaplayerui.mo
${LOC}amor.mo
${LOC}appletproxy.mo
${LOC}ark.mo
${LOC}artsbuilder.mo
${LOC}artscontrol.mo
${LOC}artsmodules.mo
${LOC}atlantik.mo
${LOC}atlantikdesigner.mo
${LOC}audiorename_plugin.mo
${LOC}autorefresh.mo
${LOC}babelfish.mo
${LOC}cervisia.mo
${LOC}charlatanui.mo
${LOC}childpanelextension.mo
${LOC}clockapplet.mo
${LOC}crashesplugin.mo
${LOC}cupsdconf.mo
${LOC}cvsservice.mo
${LOC}dcopservice.mo
${LOC}desktop_kde-i18n.mo
${LOC}desktop_kdeaccessibility.mo
${LOC}desktop_kdeaddons.mo
${LOC}desktop_kdeadmin.mo
${LOC}desktop_kdeartwork.mo
${LOC}desktop_kdebase.mo
${LOC}desktop_kdeedu.mo
${LOC}desktop_kdegames.mo
${LOC}desktop_kdegraphics.mo
${LOC}desktop_kdelibs.mo
${LOC}desktop_kdemultimedia.mo
${LOC}desktop_kdenetwork.mo
${LOC}desktop_kdepim.mo
${LOC}desktop_kdesdk.mo
${LOC}desktop_kdetoys.mo
${LOC}desktop_kdeutils.mo
${LOC}desktop_kdevelop.mo
${LOC}desktop_quanta.mo
${LOC}devicesapplet.mo
${LOC}dirfilterplugin.mo
${LOC}display.mo
${LOC}dockbarextension.mo
${LOC}domtreeviewer.mo
${LOC}drkonqi.mo
${LOC}dub.mo
${LOC}extensionproxy.mo
${LOC}ffrs.mo
${LOC}filetypes.mo
${LOC}flashkard.mo
${LOC}fontinst.mo
${LOC}fsview.mo
${LOC}htmlsearch.mo
${LOC}imagerename_plugin.mo
${LOC}imgalleryplugin.mo
${LOC}irkick.mo
${LOC}jefferson.mo
${LOC}juk.mo
${LOC}kabc2mutt.mo
${LOC}kabc_dir.mo
${LOC}kabc_file.mo
${LOC}kabc_ldap.mo
${LOC}kabc_ldapkio.mo
${LOC}kabc_net.mo
${LOC}kabc_sql.mo
${LOC}kabcformat_binary.mo
${LOC}kaboodle.mo
${LOC}kaccess.mo
${LOC}kaddressbook.mo
${LOC}kalarm.mo
${LOC}kalarmdgui.mo
${LOC}kalzium.mo
${LOC}kandy.mo
${LOC}kappfinder.mo
${LOC}karm.mo
${LOC}kasbarextension.mo
${LOC}kasteroids.mo
${LOC}kate.mo
${LOC}katecppsymbolviewer.mo
${LOC}katedefaultproject.mo
${LOC}katefll_initplugin.mo
${LOC}katefll_plugin.mo
${LOC}katehelloworld.mo
${LOC}katehtmltools.mo
${LOC}kateinsertcommand.mo
${LOC}katemake.mo
${LOC}katemodeline.mo
${LOC}kateopenheader.mo
${LOC}katepart.mo
${LOC}kateprojectmanager.mo
${LOC}katepybrowse.mo
${LOC}katespell.mo
${LOC}katetextfilter.mo
${LOC}katexmlcheck.mo
${LOC}katexmltools.mo
${LOC}katomic.mo
${LOC}kaudiocreator.mo
${LOC}kbabel.mo
${LOC}kbackgammon.mo
${LOC}kbattleship.mo
${LOC}kbinaryclock.mo
${LOC}kblackbox.mo
${LOC}kbounce.mo
${LOC}kbruch.mo
${LOC}kbugbuster.mo
${LOC}kcachegrind.mo
${LOC}kcalc.mo
${LOC}kcardchooser.mo
${LOC}kcharselect.mo
${LOC}kcharselectapplet.mo
${LOC}kcm_krfb.mo
${LOC}kcm_kviewcanvasconfig.mo
${LOC}kcm_kviewgeneralconfig.mo
${LOC}kcm_kviewpluginsconfig.mo
${LOC}kcm_kviewviewerpluginsconfig.mo
${LOC}kcmaccess.mo
${LOC}kcmaccessibility.mo
${LOC}kcmarts.mo
${LOC}kcmaudiocd.mo
${LOC}kcmbackground.mo
${LOC}kcmbell.mo
${LOC}kcmcddb.mo
${LOC}kcmcgi.mo
${LOC}kcmcolors.mo
${LOC}kcmcomponentchooser.mo
${LOC}kcmcrypto.mo
${LOC}kcmcss.mo
${LOC}kcmemail.mo
${LOC}kcmenergy.mo
${LOC}kcmfileshare.mo
${LOC}kcmfonts.mo
${LOC}kcmhtmlsearch.mo
${LOC}kcmicons.mo
${LOC}kcminfo.mo
${LOC}kcminput.mo
${LOC}kcmioslaveinfo.mo
${LOC}kcmkabconfig.mo
${LOC}kcmkamera.mo
${LOC}kcmkclock.mo
${LOC}kcmkded.mo
${LOC}kcmkeys.mo
${LOC}kcmkicker.mo
${LOC}kcmkio.mo
${LOC}kcmkmix.mo
${LOC}kcmkonq.mo
${LOC}kcmkonqhtml.mo
${LOC}kcmkonsole.mo
${LOC}kcmkontactnt.mo
${LOC}kcmktalkd.mo
${LOC}kcmkuick.mo
${LOC}kcmkurifilt.mo
${LOC}kcmkvaio.mo
${LOC}kcmkwallet.mo
${LOC}kcmkwindecoration.mo
${LOC}kcmkwintheme.mo
${LOC}kcmkwm.mo
${LOC}kcmkxmlrpcd.mo
${LOC}kcmlanbrowser.mo
${LOC}kcmlaptop.mo
${LOC}kcmlaunch.mo
${LOC}kcmlayout.mo
${LOC}kcmlilo.mo
${LOC}kcmlinuz.mo
${LOC}kcmlirc.mo
${LOC}kcmlocale.mo
${LOC}kcmmediacontrol.mo
${LOC}kcmmidi.mo
${LOC}kcmnic.mo
${LOC}kcmnotify.mo
${LOC}kcmperformance.mo
${LOC}kcmprintmgr.mo
${LOC}kcmsamba.mo
${LOC}kcmscreensaver.mo
${LOC}kcmsmartcard.mo
${LOC}kcmsmserver.mo
${LOC}kcmsocks.mo
${LOC}kcmspellchecking.mo
${LOC}kcmstyle.mo
${LOC}kcmtaskbar.mo
${LOC}kcmusb.mo
${LOC}kcmview1394.mo
${LOC}kcmvim.mo
${LOC}kcmwifi.mo
${LOC}kcmxinerama.mo
${LOC}kcoloredit.mo
${LOC}kcontrol.mo
${LOC}kcron.mo
${LOC}kdat.mo
${LOC}kdcop.mo
${LOC}kdebugdialog.mo
${LOC}kdelibs.mo
${LOC}kdelibs_colors.mo
${LOC}kdelirc.mo
${LOC}kdepasswd.mo
${LOC}kdeprint.mo
${LOC}kdeprint_part.mo
${LOC}kdeprintfax.mo
${LOC}kdesktop.mo
${LOC}kdessh.mo
${LOC}kdesu.mo
${LOC}kdesud.mo
${LOC}kdevtipofday.mo
${LOC}kdf.mo
${LOC}kdgantt.mo
${LOC}kdialog.mo
${LOC}kdict.mo
${LOC}kdictapplet.mo
${LOC}kdmchooser.mo
${LOC}kdmconfig.mo
${LOC}kdmgreet.mo
${LOC}kdvi.mo
${LOC}kedit.mo
${LOC}keduca.mo
${LOC}kenolaba.mo
${LOC}kfax.mo
${LOC}kfifteenapplet.mo
${LOC}kfile_au.mo
${LOC}kfile_avi.mo
${LOC}kfile_bmp.mo
${LOC}kfile_cpp.mo
${LOC}kfile_deb.mo
${LOC}kfile_desktop.mo
${LOC}kfile_diff.mo
${LOC}kfile_dvi.mo
${LOC}kfile_flac.mo
${LOC}kfile_folder.mo
${LOC}kfile_font.mo
${LOC}kfile_gif.mo
${LOC}kfile_html.mo
${LOC}kfile_ico.mo
${LOC}kfile_jpeg.mo
${LOC}kfile_m3u.mo
${LOC}kfile_mp3.mo
${LOC}kfile_ogg.mo
${LOC}kfile_pcx.mo
${LOC}kfile_pdf.mo
${LOC}kfile_png.mo
${LOC}kfile_pnm.mo
${LOC}kfile_po.mo
${LOC}kfile_ps.mo
${LOC}kfile_rfc822.mo
${LOC}kfile_rpm.mo
${LOC}kfile_tga.mo
${LOC}kfile_tiff.mo
${LOC}kfile_ts.mo
${LOC}kfile_txt.mo
${LOC}kfile_vcf.mo
${LOC}kfile_wav.mo
${LOC}kfile_xbm.mo
${LOC}kfileaudiopreview.mo
${LOC}kfilereplace.mo
${LOC}kfindpart.mo
${LOC}kfloppy.mo
${LOC}kfmclient.mo
${LOC}kfontinst.mo
${LOC}kfouleggs.mo
${LOC}kgamma.mo
${LOC}kgantt.mo
${LOC}kget.mo
${LOC}kghostview.mo
${LOC}kgoldrunner.mo
${LOC}kgpg.mo
${LOC}kgpgcertmanager.mo
${LOC}khangman.mo
${LOC}khelpcenter.mo
${LOC}khexedit.mo
${LOC}khotkeys.mo
${LOC}khtmlsettingsplugin.mo
${LOC}kicker.mo
${LOC}kiconedit.mo
${LOC}kig.mo
${LOC}kinetd.mo
${LOC}kio.mo
${LOC}kio_audiocd.mo
${LOC}kio_devices.mo
${LOC}kio_finger.mo
${LOC}kio_fish.mo
${LOC}kio_floppy.mo
${LOC}kio_help.mo
${LOC}kio_imap4.mo
${LOC}kio_lan.mo
${LOC}kio_mac.mo
${LOC}kio_man.mo
${LOC}kio_mobile.mo
${LOC}kio_nfs.mo
${LOC}kio_nntp.mo
${LOC}kio_pop3.mo
${LOC}kio_print.mo
${LOC}kio_settings.mo
${LOC}kio_sftp.mo
${LOC}kio_sieve.mo
${LOC}kio_smb.mo
${LOC}kio_smbro.mo
${LOC}kio_smtp.mo
${LOC}kioexec.mo
${LOC}kit.mo
${LOC}kiten.mo
${LOC}kjobviewer.mo
${LOC}kjots.mo
${LOC}kjumpingcube.mo
${LOC}klaptopdaemon.mo
${LOC}klegacyimport.mo
${LOC}klettres.mo
${LOC}klickety.mo
${LOC}klines.mo
${LOC}klipper.mo
${LOC}klock.mo
${LOC}kmag.mo
${LOC}kmahjongg.mo
${LOC}kmail.mo
${LOC}kmailcvt.mo
${LOC}kmathtool.mo
${LOC}kmcop.mo
${LOC}kmenuapplet.mo
${LOC}kmenuedit.mo
${LOC}kmessedwords.mo
${LOC}kmid.mo
${LOC}kmidi.mo
${LOC}kmines.mo
${LOC}kminipagerapplet.mo
${LOC}kmix.mo
${LOC}kmobile.mo
${LOC}kmoon.mo
${LOC}kmousetool.mo
${LOC}kmouth.mo
${LOC}kmplot.mo
${LOC}kmrml.mo
${LOC}knewsticker.mo
${LOC}knode.mo
${LOC}knorskverbs.mo
${LOC}knotes.mo
${LOC}knotify.mo
${LOC}kodo.mo
${LOC}kolf.mo
${LOC}kolourpicker.mo
${LOC}kompare.mo
${LOC}konq_smbmounterplugin.mo
${LOC}konqsidebar_mediaplayer.mo
${LOC}konqueror.mo
${LOC}konquest.mo
${LOC}konsole.mo
${LOC}konsolekalendar.mo
${LOC}kontact.mo
${LOC}kooka.mo
${LOC}kopete.mo
${LOC}korganizer.mo
${LOC}korn.mo
${LOC}kpackage.mo
${LOC}kpager.mo
${LOC}kpaint.mo
${LOC}kpartapp.mo
${LOC}kpartsaver.mo
${LOC}kpat.mo
${LOC}kpdf.mo
${LOC}kpercentage.mo
${LOC}kpersonalizer.mo
${LOC}kpf.mo
${LOC}kpilot.mo
${LOC}kpoker.mo
${LOC}kpovmodeler.mo
${LOC}kppp.mo
${LOC}kppplogview.mo
${LOC}kprinter.mo
${LOC}krandr.mo
${LOC}krdb.mo
${LOC}krdc.mo
${LOC}kreadconfig.mo
${LOC}krec.mo
${LOC}kregexpeditor.mo
${LOC}kreversi.mo
${LOC}krfb.mo
${LOC}kruler.mo
${LOC}krunapplet.mo
${LOC}ksame.mo
${LOC}kscd.mo
${LOC}kscreensaver.mo
${LOC}kshisen.mo
${LOC}ksig.mo
${LOC}ksim.mo
${LOC}ksirc.mo
${LOC}ksirtet.mo
${LOC}ksmiletris.mo
${LOC}ksmserver.mo
${LOC}ksnake.mo
${LOC}ksnapshot.mo
${LOC}ksokoban.mo
${LOC}kspaceduel.mo
${LOC}ksplash.mo
${LOC}ksplashthemes.mo
${LOC}kstars.mo
${LOC}kstart.mo
${LOC}kstartperf.mo
${LOC}kstyle_keramik_config.mo
${LOC}kstyle_plastik_config.mo
${LOC}ksvgplugin.mo
${LOC}ksync.mo
${LOC}ksysguard.mo
${LOC}ksystemtrayapplet.mo
${LOC}ksystraycmd.mo
${LOC}ksysv.mo
${LOC}ktalkd.mo
${LOC}ktaskbarapplet.mo
${LOC}kteatime.mo
${LOC}ktexteditor_insertfile.mo
${LOC}ktexteditor_isearch.mo
${LOC}ktexteditor_kdatatool.mo
${LOC}ktimemon.mo
${LOC}ktimer.mo
${LOC}ktip.mo
${LOC}ktnef.mo
${LOC}ktouch.mo
${LOC}ktron.mo
${LOC}ktuberling.mo
${LOC}ktux.mo
${LOC}kuick_plugin.mo
${LOC}kuickshow.mo
${LOC}kuiviewer.mo
${LOC}kuser.mo
${LOC}kverbos.mo
${LOC}kview.mo
${LOC}kview_scale.mo
${LOC}kviewbrowserplugin.mo
${LOC}kviewcanvas.mo
${LOC}kvieweffectsplugin.mo
${LOC}kviewpresenterplugin.mo
${LOC}kviewscannerplugin.mo
${LOC}kviewshell.mo
${LOC}kviewtemplateplugin.mo
${LOC}kviewviewer.mo
${LOC}kvoctrain.mo
${LOC}kwalletmanager.mo
${LOC}kweather.mo
${LOC}kwifimanager.mo
${LOC}kwin.mo
${LOC}kwin4.mo
${LOC}kwin_b2_config.mo
${LOC}kwin_cde_config.mo
${LOC}kwin_default_config.mo
${LOC}kwin_glow_config.mo
${LOC}kwin_icewm_config.mo
${LOC}kwin_keramik_config.mo
${LOC}kwin_modernsys_config.mo
${LOC}kwin_plastik_config.mo
${LOC}kwin_quartz_config.mo
${LOC}kwireless.mo
${LOC}kworldclock.mo
${LOC}kwriteconfig.mo
${LOC}kxkb.mo
${LOC}kxmlrpcd.mo
${LOC}kxsconfig.mo
${LOC}kxsldbg.mo
${LOC}libcalendarresources.mo
${LOC}libkaddrbk_geo_xxport.mo
${LOC}libkcal.mo
${LOC}libkcalsystem.mo
${LOC}libkcddb.mo
${LOC}libkdegames.mo
${LOC}libkdehighscores.mo
${LOC}libkdenetwork.mo
${LOC}libkdepim.mo
${LOC}libkicker.mo
${LOC}libkickermenu_kdeprint.mo
${LOC}libkickermenu_konsole.mo
${LOC}libkickermenu_prefmenu.mo
${LOC}libkickermenu_recentdocs.mo
${LOC}libkonq.mo
${LOC}libkpimexchange.mo
${LOC}libkscan.mo
${LOC}libkscreensaver.mo
${LOC}libksieve.mo
${LOC}libksirtet.mo
${LOC}libksync.mo
${LOC}libtaskbar.mo
${LOC}libtaskmanager.mo
${LOC}lockout.mo
${LOC}lskat.mo
${LOC}lyrics.mo
${LOC}mediacontrol.mo
${LOC}minitoolsplugin.mo
${LOC}naughtyapplet.mo
${LOC}nexscope.mo
${LOC}noatun.mo
${LOC}nsplugin.mo
${LOC}passwords.mo
${LOC}pitchablespeed.mo
${LOC}ppdtranslations.mo
${LOC}privacy.mo
${LOC}qeditor.mo
${LOC}quanta.mo
${LOC}quicklauncher.mo
${LOC}secpolicy.mo
${LOC}spy.mo
${LOC}synaescope.mo
${LOC}taskbarextension.mo
${LOC}timezones.mo
${LOC}tippecanoe.mo
${LOC}tyler.mo
${LOC}uachangerplugin.mo
${LOC}umbrello.mo
${LOC}userinfo.mo
${LOC}validatorsplugin.mo
${LOC}vimpart.mo
${LOC}wakeup.mo
${LOC}wavecapture.mo
${LOC}webarchiver.mo
share/locale/sv/charset
share/locale/sv/entry.desktop
share/locale/sv/flag.png
@dirrm ${DOC}umbrello/pics
@dirrm ${DOC}umbrello
@dirrm ${DOC}quanta
@dirrm ${DOC}noatun
@dirrm ${DOC}megami
@dirrm ${DOC}lskat
@dirrm ${DOC}lisa
@dirrm ${DOC}kxsldbg
@dirrm ${DOC}kxkb
@dirrm ${DOC}kxconfig
@dirrm ${DOC}kwuftpd
@dirrm ${DOC}kwrite
@dirrm ${DOC}kworldclock
@dirrm ${DOC}kwin4
@dirrm ${DOC}kwifimanager
@dirrm ${DOC}kweather
@dirrm ${DOC}kwallet
@dirrm ${DOC}kvoctrain
@dirrm ${DOC}kview
@dirrm ${DOC}kverbos
@dirrm ${DOC}kuser
@dirrm ${DOC}kuickshow
@dirrm ${DOC}ktuberling
@dirrm ${DOC}ktron
@dirrm ${DOC}ktouch
@dirrm ${DOC}ktimer
@dirrm ${DOC}kteatime
@dirrm ${DOC}ktalkd
@dirrm ${DOC}ksysv
@dirrm ${DOC}ksysguard
@dirrm ${DOC}kstars
@dirrm ${DOC}ksplashml
@dirrm ${DOC}kspell
@dirrm ${DOC}kspaceduel
@dirrm ${DOC}ksokoban
@dirrm ${DOC}ksnapshot
@dirrm ${DOC}ksnake
@dirrm ${DOC}ksirtet
@dirrm ${DOC}ksirc
@dirrm ${DOC}ksim
@dirrm ${DOC}kshisen
@dirrm ${DOC}kscd
@dirrm ${DOC}ksame
@dirrm ${DOC}kruler
@dirrm ${DOC}krfb
@dirrm ${DOC}kreversi
@dirrm ${DOC}krec
@dirrm ${DOC}krdc
@dirrm ${DOC}kppp
@dirrm ${DOC}kpovmodeler
@dirrm ${DOC}kpoker
@dirrm ${DOC}kpilot
@dirrm ${DOC}kpf
@dirrm ${DOC}kpercentage
@dirrm ${DOC}kpdf
@dirrm ${DOC}kpat
@dirrm ${DOC}kpaint
@dirrm ${DOC}kpager
@dirrm ${DOC}kpackage
@dirrm ${DOC}korn
@dirrm ${DOC}korganizer
@dirrm ${DOC}kopete
@dirrm ${DOC}kooka
@dirrm ${DOC}kontact
@dirrm ${DOC}konsolekalendar
@dirrm ${DOC}konsole
@dirrm ${DOC}konquest
@dirrm ${DOC}konqueror
@dirrm ${DOC}konq-plugins/webarchiver
@dirrm ${DOC}konq-plugins/validators
@dirrm ${DOC}konq-plugins/uachanger
@dirrm ${DOC}konq-plugins/smbmounter
@dirrm ${DOC}konq-plugins/mediaplayer
@dirrm ${DOC}konq-plugins/kuick
@dirrm ${DOC}konq-plugins/khtmlsettings
@dirrm ${DOC}konq-plugins/imgallery
@dirrm ${DOC}konq-plugins/fsview
@dirrm ${DOC}konq-plugins/domtreeviewer
@dirrm ${DOC}konq-plugins/dirfilter
@dirrm ${DOC}konq-plugins/crashes
@dirrm ${DOC}konq-plugins/babel
@dirrm ${DOC}konq-plugins
@dirrm ${DOC}kompare
@dirrm ${DOC}kolf
@dirrm ${DOC}kodo
@dirrm ${DOC}knotes
@dirrm ${DOC}knode
@dirrm ${DOC}knewsticker
@dirrm ${DOC}kmplot
@dirrm ${DOC}kmouth
@dirrm ${DOC}kmousetool
@dirrm ${DOC}kmoon
@dirrm ${DOC}kmix
@dirrm ${DOC}kmines
@dirrm ${DOC}kmidi
@dirrm ${DOC}kmid
@dirrm ${DOC}kmessedwords
@dirrm ${DOC}kmenuedit
@dirrm ${DOC}kmathtool
@dirrm ${DOC}kmail
@dirrm ${DOC}kmag/images
@dirrm ${DOC}kmag
@dirrm ${DOC}klipper
@dirrm ${DOC}klines
@dirrm ${DOC}klickety
@dirrm ${DOC}klettres
@dirrm ${DOC}kjumpingcube
@dirrm ${DOC}kjots
@dirrm ${DOC}kiten
@dirrm ${DOC}kit
@dirrm ${DOC}kioslave
@dirrm ${DOC}kinfocenter/xserver
@dirrm ${DOC}kinfocenter/usb
@dirrm ${DOC}kinfocenter/sound
@dirrm ${DOC}kinfocenter/scsi
@dirrm ${DOC}kinfocenter/samba
@dirrm ${DOC}kinfocenter/protocols
@dirrm ${DOC}kinfocenter/processor
@dirrm ${DOC}kinfocenter/pcmcia
@dirrm ${DOC}kinfocenter/pci
@dirrm ${DOC}kinfocenter/partitions
@dirrm ${DOC}kinfocenter/nics
@dirrm ${DOC}kinfocenter/memory
@dirrm ${DOC}kinfocenter/ioports
@dirrm ${DOC}kinfocenter/interrupts
@dirrm ${DOC}kinfocenter/dma
@dirrm ${DOC}kinfocenter/devices
@dirrm ${DOC}kinfocenter/blockdevices
@dirrm ${DOC}kinfocenter
@dirrm ${DOC}kig
@dirrm ${DOC}kiconedit
@dirrm ${DOC}kicker-applets
@dirrm ${DOC}kicker
@dirrm ${DOC}khexedit
@dirrm ${DOC}khelpcenter/visualdict
@dirrm ${DOC}khelpcenter/userguide
@dirrm ${DOC}khelpcenter/quickstart
@dirrm ${DOC}khelpcenter/glossary
@dirrm ${DOC}khelpcenter/faq
@dirrm ${DOC}khelpcenter
@dirrm ${DOC}khangman
@dirrm ${DOC}kgpgcertmanager
@dirrm ${DOC}kgpg
@dirrm ${DOC}kgoldrunner
@dirrm ${DOC}kghostview
@dirrm ${DOC}kget
@dirrm ${DOC}kgamma
@dirrm ${DOC}kfouleggs
@dirrm ${DOC}kfloppy
@dirrm ${DOC}kfind
@dirrm ${DOC}kenolaba
@dirrm ${DOC}keduca
@dirrm ${DOC}kedit
@dirrm ${DOC}kdvi
@dirrm ${DOC}kdm
@dirrm ${DOC}kdict
@dirrm ${DOC}kdf
@dirrm ${DOC}kdesu
@dirrm ${DOC}kdeprint
@dirrm ${DOC}kdebugdialog
@dirrm ${DOC}kdat
@dirrm ${DOC}kcron
@dirrm ${DOC}kcontrol/windowmanagement
@dirrm ${DOC}kcontrol/useragent
@dirrm ${DOC}kcontrol/spellchecking
@dirrm ${DOC}kcontrol/smb
@dirrm ${DOC}kcontrol/screensaver
@dirrm ${DOC}kcontrol/proxy
@dirrm ${DOC}kcontrol/powerctrl
@dirrm ${DOC}kcontrol/passwords
@dirrm ${DOC}kcontrol/panelappearance
@dirrm ${DOC}kcontrol/panel
@dirrm ${DOC}kcontrol/netpref
@dirrm ${DOC}kcontrol/mouse
@dirrm ${DOC}kcontrol/laptop
@dirrm ${DOC}kcontrol/language
@dirrm ${DOC}kcontrol/lanbrowser
@dirrm ${DOC}kcontrol/kxmlrpcd
@dirrm ${DOC}kcontrol/kwindecoration
@dirrm ${DOC}kcontrol/kthememgr
@dirrm ${DOC}kcontrol/kmixcfg
@dirrm ${DOC}kcontrol/khtml
@dirrm ${DOC}kcontrol/keys
@dirrm ${DOC}kcontrol/keyboard
@dirrm ${DOC}kcontrol/kdm
@dirrm ${DOC}kcontrol/kcmtaskbar
@dirrm ${DOC}kcontrol/kcmstyle
@dirrm ${DOC}kcontrol/kcmsmserver
@dirrm ${DOC}kcontrol/kcmnotify
@dirrm ${DOC}kcontrol/kcmlowbatwarn
@dirrm ${DOC}kcontrol/kcmlowbatcrit
@dirrm ${DOC}kcontrol/kcmlaunch
@dirrm ${DOC}kcontrol/kcmktalkd
@dirrm ${DOC}kcontrol/kcmkonsole
@dirrm ${DOC}kcontrol/kcmfontinst
@dirrm ${DOC}kcontrol/kcmcss
@dirrm ${DOC}kcontrol/kcmaccess
@dirrm ${DOC}kcontrol/kalarmd
@dirrm ${DOC}kcontrol/icons
@dirrm ${DOC}kcontrol/helpindex
@dirrm ${DOC}kcontrol/fonts
@dirrm ${DOC}kcontrol/filetypes
@dirrm ${DOC}kcontrol/filemanager
@dirrm ${DOC}kcontrol/energy
@dirrm ${DOC}kcontrol/email
@dirrm ${DOC}kcontrol/ebrowsing
@dirrm ${DOC}kcontrol/desktopbehavior
@dirrm ${DOC}kcontrol/desktop
@dirrm ${DOC}kcontrol/crypto
@dirrm ${DOC}kcontrol/cookies
@dirrm ${DOC}kcontrol/colors
@dirrm ${DOC}kcontrol/clock
@dirrm ${DOC}kcontrol/cache
@dirrm ${DOC}kcontrol/bell
@dirrm ${DOC}kcontrol/background
@dirrm ${DOC}kcontrol/arts
@dirrm ${DOC}kcontrol
@dirrm ${DOC}kcoloredit
@dirrm ${DOC}kcharselect
@dirrm ${DOC}kcalc
@dirrm ${DOC}kcachegrind
@dirrm ${DOC}kbugbuster
@dirrm ${DOC}kbruch
@dirrm ${DOC}kbounce
@dirrm ${DOC}kblackbox
@dirrm ${DOC}kbattleship
@dirrm ${DOC}kbackgammon
@dirrm ${DOC}kbabel
@dirrm ${DOC}katomic
@dirrm ${DOC}kate-plugins
@dirrm ${DOC}kate
@dirrm ${DOC}kasteroids
@dirrm ${DOC}karm
@dirrm ${DOC}kandy
@dirrm ${DOC}kamera
@dirrm ${DOC}kalzium
@dirrm ${DOC}kalarm
@dirrm ${DOC}kaddressbook
@dirrm ${DOC}kaboodle
@dirrm ${DOC}juk
@dirrm ${DOC}flashkard
@dirrm ${DOC}common
@dirrm ${DOC}cervisia
@dirrm ${DOC}atlantik
@dirrm ${DOC}artsbuilder/images
@dirrm ${DOC}artsbuilder
@dirrm ${DOC}ark
@dirrm ${DOC}amor
@dirrm ${DOC}KRegExpEditor
@dirrm share/doc/HTML/sv
@dirrm share/apps/ktuberling/sounds/sv
@dirrm share/apps/ktuberling/sounds
@dirrm share/apps/ktuberling
